.subckt vddtie vdd vss z
*04-JAN-08 SPICE3       file   created      from vddtie.ext -        technology: scmos
m00 z vss vdd vdd p w=1.65u  l=0.13u ad=0.80025p  pd=4.27u as=0.80025p  ps=4.27u
m01 z vss vss vss n w=1.265u l=0.13u ad=0.613525p pd=3.5u  as=0.613525p ps=3.5u 
C0  z   w1  0.013f
C1  vdd w2  0.030f
C2  z   w3  0.022f
C3  z   w4  0.010f
C4  z   w2  0.030f
C5  w1  w2  0.166f
C6  w3  w2  0.166f
C7  w4  w2  0.166f
C8  vdd z   0.057f
C9  vdd w1  0.013f
C10 vdd w3  0.005f
C11 w2  vss 1.078f
C12 w4  vss 0.200f
C13 w3  vss 0.185f
C14 w1  vss 0.186f
C15 z   vss 0.107f
.ends
