.subckt o3_x4 i0 i1 i2 q vdd vss
*05-JAN-08 SPICE3       file   created      from o3_x4.ext -        technology: scmos
m00 w1  i2 w2  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.697p    ps=4.13u   
m01 w3  i1 w1  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.2542p   ps=1.95u   
m02 vdd i0 w3  vdd p w=1.64u l=0.13u ad=0.750913p pd=3.08658u as=0.2542p   ps=1.95u   
m03 q   w2 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=1.00274p  ps=4.12171u
m04 vdd w2 q   vdd p w=2.19u l=0.13u ad=1.00274p  pd=4.12171u as=0.58035p  ps=2.72u   
m05 vss i2 w2  vss n w=0.54u l=0.13u ad=0.191643p pd=1.35142u as=0.1719p   ps=1.35667u
m06 w2  i1 vss vss n w=0.54u l=0.13u ad=0.1719p   pd=1.35667u as=0.191643p ps=1.35142u
m07 vss i0 w2  vss n w=0.54u l=0.13u ad=0.191643p pd=1.35142u as=0.1719p   ps=1.35667u
m08 q   w2 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.386835p ps=2.72787u
m09 vss w2 q   vss n w=1.09u l=0.13u ad=0.386835p pd=2.72787u as=0.28885p  ps=1.62u   
C0  w2  i2  0.048f
C1  vdd i0  0.022f
C2  w2  i1  0.028f
C3  w2  i0  0.178f
C4  i2  i1  0.240f
C5  w2  w1  0.008f
C6  vdd q   0.076f
C7  w2  w3  0.008f
C8  i1  i0  0.223f
C9  w2  q   0.159f
C10 i1  w1  0.012f
C11 i1  w3  0.012f
C12 vdd w2  0.155f
C13 vdd i2  0.002f
C14 vdd i1  0.002f
C15 q   vss 0.144f
C16 w3  vss 0.010f
C17 w1  vss 0.010f
C18 i0  vss 0.130f
C19 i1  vss 0.119f
C20 i2  vss 0.126f
C21 w2  vss 0.430f
.ends
