.subckt aoi21bv0x05 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from aoi21bv0x05.ext -        technology: scmos
m00 n1  bn z   vdd p w=0.88u  l=0.13u ad=0.213033p  pd=1.70333u  as=0.31185p   ps=2.51u    
m01 vdd a2 n1  vdd p w=0.88u  l=0.13u ad=0.3806p    pd=2.89818u  as=0.213033p  ps=1.70333u 
m02 n1  a1 vdd vdd p w=0.88u  l=0.13u ad=0.213033p  pd=1.70333u  as=0.3806p    ps=2.89818u 
m03 vdd b  bn  vdd p w=0.66u  l=0.13u ad=0.28545p   pd=2.17364u  as=0.2112p    ps=2.07u    
m04 z   bn vss vss n w=0.33u  l=0.13u ad=0.0706962p pd=0.743077u as=0.136168p  ps=1.23158u 
m05 w1  a2 z   vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u     as=0.0824789p ps=0.866923u
m06 vss a1 w1  vss n w=0.385u l=0.13u ad=0.158863p  pd=1.43684u  as=0.0490875p ps=0.64u    
m07 bn  b  vss vss n w=0.33u  l=0.13u ad=0.12375p   pd=1.41u     as=0.136168p  ps=1.23158u 
C0  vdd n1  0.088f
C1  a1  a2  0.118f
C2  a1  z   0.006f
C3  vdd b   0.034f
C4  bn  a2  0.204f
C5  bn  z   0.062f
C6  a1  n1  0.030f
C7  a2  z   0.047f
C8  a1  b   0.023f
C9  bn  b   0.093f
C10 a2  n1  0.007f
C11 z   n1  0.007f
C12 a2  w1  0.007f
C13 vdd a1  0.023f
C14 a1  bn  0.093f
C15 w1  vss 0.001f
C16 b   vss 0.120f
C17 n1  vss 0.037f
C18 z   vss 0.224f
C19 a2  vss 0.156f
C20 bn  vss 0.170f
C21 a1  vss 0.102f
.ends
