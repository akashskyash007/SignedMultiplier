.subckt cgi2bv0x3 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from cgi2bv0x3.ext -        technology: scmos
m00 vdd b  bn  vdd p w=0.44u l=0.13u ad=0.108329p pd=0.612152u as=0.0999625p ps=0.69375u
m01 bn  b  vdd vdd p w=1.54u l=0.13u ad=0.349869p pd=2.42813u  as=0.379152p  ps=2.14253u
m02 vdd b  bn  vdd p w=1.54u l=0.13u ad=0.379152p pd=2.14253u  as=0.349869p  ps=2.42813u
m03 n1  bn vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u  as=0.379152p  ps=2.14253u
m04 vdd bn n1  vdd p w=1.54u l=0.13u ad=0.379152p pd=2.14253u  as=0.34155p   ps=2.16778u
m05 n1  bn vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u  as=0.379152p  ps=2.14253u
m06 z   c  n1  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u     as=0.34155p   ps=2.16778u
m07 n1  c  z   vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u  as=0.3234p    ps=1.96u   
m08 z   c  n1  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u     as=0.34155p   ps=2.16778u
m09 w1  bn z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u    as=0.3234p    ps=1.96u   
m10 vdd a  w1  vdd p w=1.54u l=0.13u ad=0.379152p pd=2.14253u  as=0.19635p   ps=1.795u  
m11 w2  a  vdd vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u    as=0.379152p  ps=2.14253u
m12 z   bn w2  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u     as=0.19635p   ps=1.795u  
m13 w3  bn z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u    as=0.3234p    ps=1.96u   
m14 vdd a  w3  vdd p w=1.54u l=0.13u ad=0.379152p pd=2.14253u  as=0.19635p   ps=1.795u  
m15 n1  a  vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u  as=0.379152p  ps=2.14253u
m16 vdd a  n1  vdd p w=1.54u l=0.13u ad=0.379152p pd=2.14253u  as=0.34155p   ps=2.16778u
m17 n1  a  vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u  as=0.379152p  ps=2.14253u
m18 bn  b  vss vss n w=0.88u l=0.13u ad=0.1848p   pd=1.3u      as=0.280669p  ps=1.80718u
m19 vss b  bn  vss n w=0.88u l=0.13u ad=0.280669p pd=1.80718u  as=0.1848p    ps=1.3u    
m20 n3  bn vss vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u  as=0.245586p  ps=1.58128u
m21 vss bn n3  vss n w=0.77u l=0.13u ad=0.245586p pd=1.58128u  as=0.1617p    ps=1.14935u
m22 n3  bn vss vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u  as=0.245586p  ps=1.58128u
m23 z   c  n3  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u     as=0.1617p    ps=1.14935u
m24 n3  c  z   vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u  as=0.1617p    ps=1.19u   
m25 z   c  n3  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u     as=0.1617p    ps=1.14935u
m26 w4  bn z   vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u    as=0.1617p    ps=1.19u   
m27 vss a  w4  vss n w=0.77u l=0.13u ad=0.245586p pd=1.58128u  as=0.098175p  ps=1.025u  
m28 w5  a  vss vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u    as=0.245586p  ps=1.58128u
m29 z   bn w5  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u     as=0.098175p  ps=1.025u  
m30 w6  bn z   vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u    as=0.1617p    ps=1.19u   
m31 vss a  w6  vss n w=0.77u l=0.13u ad=0.245586p pd=1.58128u  as=0.098175p  ps=1.025u  
m32 n3  a  vss vss n w=1.1u  l=0.13u ad=0.231p    pd=1.64194u  as=0.350837p  ps=2.25897u
m33 vss a  n3  vss n w=1.1u  l=0.13u ad=0.350837p pd=2.25897u  as=0.231p     ps=1.64194u
C0  w3  a   0.006f
C1  n3  bn  0.136f
C2  bn  z   0.073f
C3  c   n1  0.044f
C4  w3  n1  0.008f
C5  n3  c   0.044f
C6  w4  bn  0.007f
C7  c   z   0.117f
C8  a   n1  0.037f
C9  w3  z   0.009f
C10 n3  a   0.030f
C11 w5  bn  0.007f
C12 a   z   0.291f
C13 vdd b   0.019f
C14 n1  z   0.395f
C15 w2  a   0.006f
C16 vdd bn  0.101f
C17 n3  z   0.334f
C18 n1  w1  0.008f
C19 w2  n1  0.008f
C20 vdd c   0.021f
C21 n3  w4  0.008f
C22 z   w1  0.009f
C23 w2  z   0.009f
C24 w3  vdd 0.004f
C25 vdd a   0.061f
C26 b   bn  0.202f
C27 n3  w5  0.008f
C28 vdd n1  0.478f
C29 n3  w6  0.008f
C30 w6  z   0.009f
C31 vdd z   0.081f
C32 bn  c   0.185f
C33 vdd w1  0.004f
C34 bn  a   0.504f
C35 w2  vdd 0.004f
C36 bn  n1  0.031f
C37 w6  vss 0.003f
C38 w5  vss 0.004f
C39 w4  vss 0.004f
C40 n3  vss 0.538f
C41 w3  vss 0.006f
C42 w2  vss 0.007f
C43 w1  vss 0.007f
C44 z   vss 0.221f
C45 n1  vss 0.158f
C46 a   vss 0.388f
C47 c   vss 0.199f
C48 bn  vss 0.699f
C49 b   vss 0.274f
.ends
