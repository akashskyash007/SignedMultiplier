.subckt nr2a_x05 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2a_x05.ext -        technology: scmos
m00 w1  b  z   vdd p w=1.21u  l=0.13u ad=0.18755p  pd=1.52u    as=0.4477p   ps=3.28u   
m01 vdd an w1  vdd p w=1.21u  l=0.13u ad=0.421328p pd=2.08718u as=0.18755p  ps=1.52u   
m02 an  a  vdd vdd p w=0.935u l=0.13u ad=0.374825p pd=2.73u    as=0.325572p ps=1.61282u
m03 z   b  vss vss n w=0.33u  l=0.13u ad=0.08745p  pd=0.86u    as=0.173879p ps=1.36571u
m04 vss an z   vss n w=0.33u  l=0.13u ad=0.173879p pd=1.36571u as=0.08745p  ps=0.86u   
m05 an  a  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.260818p ps=2.04857u
C0  vdd w2  0.038f
C1  b   w3  0.002f
C2  an  w4  0.002f
C3  z   a   0.041f
C4  z   w4  0.001f
C5  b   w5  0.015f
C6  an  w3  0.012f
C7  w1  a   0.033f
C8  b   w2  0.014f
C9  w1  w4  0.001f
C10 an  w5  0.033f
C11 z   w3  0.012f
C12 an  w2  0.023f
C13 z   w5  0.009f
C14 vdd an  0.005f
C15 z   w2  0.053f
C16 a   w3  0.033f
C17 w1  w2  0.002f
C18 b   an  0.160f
C19 a   w2  0.019f
C20 b   z   0.099f
C21 vdd a   0.049f
C22 w4  w2  0.166f
C23 vdd w4  0.010f
C24 w3  w2  0.166f
C25 vdd w3  0.004f
C26 b   a   0.031f
C27 w5  w2  0.166f
C28 b   w4  0.002f
C29 an  a   0.145f
C30 w2  vss 1.030f
C31 w5  vss 0.177f
C32 w3  vss 0.172f
C33 w4  vss 0.188f
C34 a   vss 0.081f
C35 z   vss 0.106f
C36 an  vss 0.130f
C37 b   vss 0.123f
.ends
