* Spice description of aoi22_x1
* Spice driver version 134999461
* Date  4/01/2008 at 18:51:14
* vxlib 0.13um values
.subckt aoi22_x1 a1 a2 b1 b2 vdd vss z
M1  sig5  b1    z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2  vdd   a1    sig5  vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3  z     b2    sig5  vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M4  sig5  a2    vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M5  n2    b1    vss   vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M6  vss   a1    sig3  vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M7  z     b2    n2    vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M8  sig3  a2    z     vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
C9  a1    vss   0.789f
C8  a2    vss   0.756f
C7  b1    vss   0.742f
C10 b2    vss   0.789f
C5  sig5  vss   0.521f
C4  z     vss   1.032f
.ends
