.subckt bf1v6x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v6x2.ext -        technology: scmos
m00 vdd an z   vdd p w=1.485u l=0.13u ad=0.493763p pd=2.74295u as=0.472175p ps=3.72u   
m01 an  a  vdd vdd p w=0.935u l=0.13u ad=0.284075p pd=2.62u    as=0.310888p ps=1.72705u
m02 vss an z   vss n w=0.66u  l=0.13u ad=0.21846p  pd=1.56u    as=0.2112p   ps=2.07u   
m03 an  a  vss vss n w=0.44u  l=0.13u ad=0.1529p   pd=1.63u    as=0.14564p  ps=1.04u   
C0 vdd an  0.031f
C1 vdd z   0.049f
C2 an  z   0.133f
C3 an  a   0.151f
C4 a   vss 0.100f
C5 z   vss 0.196f
C6 an  vss 0.143f
.ends
