.subckt oai21v0x1 a1 a2 b vdd vss z
*10-JAN-08 SPICE3       file   created      from oai21v0x1.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.43u l=0.13u ad=0.431383p pd=2.51u    as=0.53625p  ps=3.61u   
m01 w2  a1  vdd vdd p w=1.43u l=0.13u ad=0.53625p  pd=3.61u    as=0.431383p ps=2.51u   
m02 z   a2  w2  vdd p w=1.43u l=0.13u ad=0.37895p  pd=1.96u    as=0.53625p  ps=3.61u   
m03 vdd b   z   vdd p w=1.43u l=0.13u ad=0.431383p pd=2.51u    as=0.37895p  ps=1.96u   
m04 vss vss w3  vss n w=0.99u l=0.13u ad=0.29865p  pd=1.92333u as=0.37125p  ps=2.73u   
m05 w4  a1  vss vss n w=0.99u l=0.13u ad=0.29865p  pd=1.92333u as=0.29865p  ps=1.92333u
m06 w4  a2  vss vss n w=0.99u l=0.13u ad=0.29865p  pd=1.92333u as=0.29865p  ps=1.92333u
m07 z   b   w4  vss n w=0.99u l=0.13u ad=0.37125p  pd=2.73u    as=0.29865p  ps=1.92333u
C0  vdd b   0.031f
C1  a1  a2  0.046f
C2  z   w4  0.041f
C3  vdd w2  0.043f
C4  vdd z   0.009f
C5  a2  b   0.129f
C6  a1  w2  0.017f
C7  a2  w2  0.001f
C8  a2  z   0.098f
C9  b   z   0.152f
C10 a2  w4  0.006f
C11 vdd a1  0.100f
C12 w2  z   0.009f
C13 vdd a2  0.009f
C14 w4  vss 0.168f
C15 w3  vss 0.011f
C16 z   vss 0.088f
C17 w2  vss 0.052f
C18 w1  vss 0.014f
C19 b   vss 0.193f
C20 a2  vss 0.207f
C21 a1  vss 0.302f
.ends
