* Spice description of xnr2_x05
* Spice driver version 134999461
* Date  4/01/2008 at 19:17:39
* vxlib 0.13um values
.subckt xnr2_x05 a b vdd vss z
M1  vdd   sig3  1     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2  1     sig4  z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M3  z     b     sig3  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M4  sig3  a     vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M5  vdd   b     sig4  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M6  z     sig3  sig4  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M7  sig3  sig4  z     vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M8  vss   a     sig3  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M9  sig4  b     vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
C5  a     vss   0.860f
C6  b     vss   1.036f
C3  sig3  vss   0.977f
C4  sig4  vss   1.455f
C2  z     vss   0.972f
.ends
