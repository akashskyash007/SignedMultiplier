* Spice description of nr2_x05
* Spice driver version 134999461
* Date  4/01/2008 at 19:07:31
* vsxlib 0.13um values
.subckt nr2_x05 a b vdd vss z
M1  n1    b     z     vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M2  vdd   a     n1    vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M3  vss   b     z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M4  z     a     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C4  a     vss   0.669f
C3  b     vss   0.833f
C2  z     vss   0.644f
.ends
