.subckt bf1v5x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v5x2.ext -        technology: scmos
m00 vdd an z   vdd p w=1.54u l=0.13u ad=0.3234p  pd=1.96u as=0.48675p ps=3.83u
m01 an  a  vdd vdd p w=1.54u l=0.13u ad=0.4444p  pd=3.83u as=0.3234p  ps=1.96u
m02 vss an z   vss n w=0.77u l=0.13u ad=0.1617p  pd=1.19u as=0.28875p ps=2.29u
m03 an  a  vss vss n w=0.77u l=0.13u ad=0.28875p pd=2.29u as=0.1617p  ps=1.19u
C0 an a   0.180f
C1 an z   0.141f
C2 an vdd 0.039f
C3 a  vdd 0.007f
C4 z  vdd 0.056f
C6 z  vss 0.196f
C7 a  vss 0.102f
C8 an vss 0.174f
.ends
