* Spice description of bf1_x1
* Spice driver version 134999461
* Date  4/01/2008 at 18:53:35
* vsxlib 0.13um values
.subckt bf1_x1 a vdd vss z
M1a 2z    a     vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M1z vdd   2z    z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2a vss   a     2z    vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M2z z     2z    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C3  2z    vss   0.954f
C4  a     vss   0.681f
C1  z     vss   0.506f
.ends
