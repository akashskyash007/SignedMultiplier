* Spice description of oa2ao222_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:33:53
* sxlib 0.13um values
.subckt oa2ao222_x2 i0 i1 i2 i3 i4 q vdd vss
Mtr_00001 vss   sig2  q     vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 vss   i2    sig1  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00003 sig1  i3    vss   vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00004 sig2  i1    sig4  vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00005 sig4  i0    vss   vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00006 sig1  i4    sig2  vss n  L=0.12U  W=0.65U  AS=0.17225P  AD=0.17225P  PS=1.83U   PD=1.83U
Mtr_00007 q     sig2  vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00008 sig6  i3    sig5  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00009 sig6  i1    vdd   vdd p  L=0.12U  W=1.585U AS=0.420025P AD=0.420025P PS=3.7U    PD=3.7U
Mtr_00010 vdd   i0    sig6  vdd p  L=0.12U  W=1.585U AS=0.420025P AD=0.420025P PS=3.7U    PD=3.7U
Mtr_00011 sig5  i2    sig2  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00012 sig2  i4    sig6  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C8  i0    vss   0.766f
C12 i1    vss   0.699f
C9  i2    vss   0.598f
C11 i3    vss   0.563f
C10 i4    vss   0.654f
C13 q     vss   0.811f
C1  sig1  vss   0.182f
C2  sig2  vss   1.019f
C6  sig6  vss   0.369f
.ends
