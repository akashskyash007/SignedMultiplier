.subckt aoi22_x1 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from aoi22_x1.ext -        technology: scmos
m00 z   b1 n3  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u  as=0.6138p   ps=3.9125u
m01 n3  b2 z   vdd p w=2.145u l=0.13u ad=0.6138p   pd=3.9125u as=0.568425p ps=2.675u 
m02 vdd a2 n3  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u  as=0.6138p   ps=3.9125u
m03 n3  a1 vdd vdd p w=2.145u l=0.13u ad=0.6138p   pd=3.9125u as=0.568425p ps=2.675u 
m04 w1  b1 vss vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u  as=0.518513p ps=3.335u 
m05 z   b2 w1  vss n w=0.935u l=0.13u ad=0.247775p pd=1.465u  as=0.144925p ps=1.245u 
m06 w2  a2 z   vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u  as=0.247775p ps=1.465u 
m07 vss a1 w2  vss n w=0.935u l=0.13u ad=0.518513p pd=3.335u  as=0.144925p ps=1.245u 
C0  b2 z   0.060f
C1  b1 vdd 0.010f
C2  z  w1  0.009f
C3  b1 b2  0.187f
C4  b1 w1  0.012f
C5  b2 vdd 0.010f
C6  a2 vdd 0.034f
C7  b1 a1  0.019f
C8  b2 a2  0.165f
C9  n3 z   0.105f
C10 a1 vdd 0.010f
C11 b1 n3  0.007f
C12 b2 a1  0.003f
C13 n3 vdd 0.177f
C14 b2 n3  0.042f
C15 a2 a1  0.202f
C16 a1 w2  0.012f
C17 a2 n3  0.064f
C18 a1 n3  0.007f
C19 b1 z   0.183f
C20 z  vdd 0.017f
C21 w2 vss 0.006f
C22 w1 vss 0.002f
C24 z  vss 0.242f
C25 n3 vss 0.100f
C26 a1 vss 0.128f
C27 a2 vss 0.120f
C28 b2 vss 0.127f
C29 b1 vss 0.115f
.ends
