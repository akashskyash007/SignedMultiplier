.subckt xaon22_x1 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon22_x1.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.925u l=0.13u ad=0.721875p pd=2.675u   as=0.552475p ps=3.20667u
m01 an  a2 vdd vdd p w=1.925u l=0.13u ad=0.552475p pd=3.20667u as=0.721875p ps=2.675u  
m02 z   bn an  vdd p w=1.925u l=0.13u ad=0.510125p pd=2.455u   as=0.552475p ps=3.20667u
m03 bn  an z   vdd p w=1.925u l=0.13u ad=0.693642p pd=3.35333u as=0.510125p ps=2.455u  
m04 vdd b1 bn  vdd p w=1.925u l=0.13u ad=0.721875p pd=2.675u   as=0.693642p ps=3.35333u
m05 bn  b2 vdd vdd p w=1.925u l=0.13u ad=0.693642p pd=3.35333u as=0.721875p ps=2.675u  
m06 w1  a1 vss vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.679276p ps=3.6523u 
m07 an  a2 w1  vss n w=1.815u l=0.13u ad=0.480975p pd=2.76375u as=0.281325p ps=2.125u  
m08 w2  b2 an  vss n w=1.265u l=0.13u ad=0.196075p pd=1.575u   as=0.335225p ps=1.92625u
m09 z   b1 w2  vss n w=1.265u l=0.13u ad=0.335225p pd=2.0139u  as=0.196075p ps=1.575u  
m10 w3  bn z   vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.26235p  ps=1.5761u 
m11 vss an w3  vss n w=0.99u  l=0.13u ad=0.370514p pd=1.99216u as=0.15345p  ps=1.3u    
m12 w4  b1 vss vss n w=1.265u l=0.13u ad=0.196075p pd=1.575u   as=0.473435p ps=2.54554u
m13 bn  b2 w4  vss n w=1.265u l=0.13u ad=0.389675p pd=3.39u    as=0.196075p ps=1.575u  
C0  vdd a1  0.010f
C1  b2  a2  0.028f
C2  an  b1  0.046f
C3  w5  w6  0.166f
C4  b2  w6  0.049f
C5  z   w7  0.012f
C6  w6  a2  0.017f
C7  w5  bn  0.009f
C8  b2  vdd 0.010f
C9  vdd a2  0.024f
C10 b2  bn  0.048f
C11 a2  bn  0.057f
C12 b1  w8  0.001f
C13 vdd w6  0.064f
C14 z   w5  0.009f
C15 an  w2  0.010f
C16 w6  bn  0.038f
C17 b2  z   0.016f
C18 z   a2  0.067f
C19 vdd bn  0.169f
C20 b1  w7  0.015f
C21 an  w3  0.020f
C22 z   w6  0.037f
C23 vdd z   0.017f
C24 z   bn  0.029f
C25 b1  w5  0.002f
C26 w1  w5  0.002f
C27 b1  b2  0.278f
C28 b1  w6  0.027f
C29 an  w8  0.046f
C30 b1  vdd 0.060f
C31 w1  w6  0.009f
C32 b1  bn  0.168f
C33 w2  w6  0.004f
C34 an  w7  0.020f
C35 b1  z   0.008f
C36 an  a1  0.007f
C37 w3  w6  0.003f
C38 an  w5  0.029f
C39 b2  w4  0.026f
C40 z   w2  0.015f
C41 an  b2  0.016f
C42 an  a2  0.092f
C43 w8  a1  0.002f
C44 w4  w6  0.002f
C45 an  w6  0.101f
C46 b2  w8  0.001f
C47 an  vdd 0.180f
C48 w7  a1  0.002f
C49 w8  a2  0.001f
C50 an  bn  0.349f
C51 w8  w6  0.166f
C52 b2  w7  0.002f
C53 vdd w8  0.022f
C54 an  z   0.294f
C55 w5  a1  0.011f
C56 w7  a2  0.030f
C57 w8  bn  0.046f
C58 a1  a2  0.161f
C59 w7  w6  0.166f
C60 z   w8  0.005f
C61 b2  w5  0.019f
C62 vdd w7  0.006f
C63 w6  a1  0.019f
C64 w5  a2  0.012f
C65 w7  bn  0.025f
C66 w6  vss 0.916f
C67 w5  vss 0.166f
C68 w7  vss 0.154f
C69 w8  vss 0.143f
C70 w1  vss 0.010f
C71 z   vss 0.017f
C73 b2  vss 0.323f
C74 b1  vss 0.169f
C75 an  vss 0.205f
C76 bn  vss 0.133f
C77 a2  vss 0.082f
C78 a1  vss 0.111f
.ends
