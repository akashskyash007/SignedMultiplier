.subckt vfeed2 vdd vss
*01-JAN-08 SPICE3       file   created      from vfeed2.ext -        technology: scmos
.ends
