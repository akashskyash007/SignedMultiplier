.subckt aoi21v0x1 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from aoi21v0x1.ext -        technology: scmos
m00 n1  b  z   vdd p w=1.485u l=0.13u ad=0.365292p  pd=2.51u    as=0.472175p ps=3.72u   
m01 vdd a2 n1  vdd p w=1.485u l=0.13u ad=0.31185p   pd=1.905u   as=0.365292p ps=2.51u   
m02 n1  a1 vdd vdd p w=1.485u l=0.13u ad=0.365292p  pd=2.51u    as=0.31185p  ps=1.905u  
m03 z   b  vss vss n w=0.385u l=0.13u ad=0.0864224p pd=0.79579u as=0.255822p ps=1.89u   
m04 w1  a2 z   vss n w=0.66u  l=0.13u ad=0.08415p   pd=0.915u   as=0.148153p ps=1.36421u
m05 vss a1 w1  vss n w=0.66u  l=0.13u ad=0.438553p  pd=3.24u    as=0.08415p  ps=0.915u  
C0  b  z   0.068f
C1  a2 a1  0.172f
C2  b  n1  0.058f
C3  a2 z   0.008f
C4  b  vdd 0.014f
C5  a1 z   0.007f
C6  a2 n1  0.025f
C7  a1 n1  0.006f
C8  a2 vdd 0.007f
C9  z  n1  0.036f
C10 a1 vdd 0.007f
C11 z  vdd 0.022f
C12 n1 vdd 0.097f
C13 b  a2  0.126f
C14 z  w1  0.004f
C15 w1 vss 0.007f
C17 n1 vss 0.049f
C18 z  vss 0.282f
C19 a1 vss 0.123f
C20 a2 vss 0.115f
C21 b  vss 0.090f
.ends
