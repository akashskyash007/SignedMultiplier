.subckt aon21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from aon21_x1.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.1u   l=0.13u ad=0.341917p pd=2.06111u  as=0.34595p  ps=3.06u   
m01 n2  b  zn  vdd p w=1.43u  l=0.13u ad=0.3971p   pd=2.54667u  as=0.4334p   ps=3.72u   
m02 vdd a2 n2  vdd p w=1.43u  l=0.13u ad=0.444492p pd=2.67944u  as=0.3971p   ps=2.54667u
m03 n2  a1 vdd vdd p w=1.43u  l=0.13u ad=0.3971p   pd=2.54667u  as=0.444492p ps=2.67944u
m04 vss zn z   vss n w=0.55u  l=0.13u ad=0.267793p pd=1.76207u  as=0.2002p   ps=1.96u   
m05 zn  b  vss vss n w=0.385u l=0.13u ad=0.102025p pd=0.876842u as=0.187455p ps=1.23345u
m06 w1  a2 zn  vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u     as=0.1749p   ps=1.50316u
m07 vss a1 w1  vss n w=0.66u  l=0.13u ad=0.321352p pd=2.11448u  as=0.1023p   ps=0.97u   
C0  w2  z   0.009f
C1  zn  w3  0.010f
C2  z   w4  0.004f
C3  vdd zn  0.006f
C4  w2  w5  0.166f
C5  w5  w4  0.166f
C6  z   w3  0.009f
C7  n2  w4  0.035f
C8  a1  w1  0.014f
C9  vdd z   0.029f
C10 b   a2  0.157f
C11 w5  w3  0.166f
C12 w2  a1  0.024f
C13 w5  vdd 0.046f
C14 a1  w4  0.001f
C15 vdd n2  0.106f
C16 b   zn  0.085f
C17 vdd a1  0.007f
C18 w5  b   0.015f
C19 b   n2  0.070f
C20 w5  a2  0.013f
C21 vdd w4  0.016f
C22 zn  z   0.052f
C23 a2  n2  0.031f
C24 w5  zn  0.031f
C25 a2  a1  0.190f
C26 w5  z   0.027f
C27 w2  b   0.001f
C28 b   w4  0.002f
C29 zn  a1  0.034f
C30 w5  n2  0.007f
C31 w2  a2  0.002f
C32 a2  w4  0.001f
C33 b   w3  0.011f
C34 vdd b   0.022f
C35 w5  a1  0.031f
C36 w2  zn  0.022f
C37 a2  w3  0.033f
C38 zn  w4  0.006f
C39 n2  a1  0.007f
C40 vdd a2  0.012f
C41 w5  vss 1.020f
C42 w2  vss 0.177f
C43 w3  vss 0.177f
C44 w4  vss 0.164f
C45 a1  vss 0.163f
C46 n2  vss 0.001f
C47 z   vss 0.042f
C48 zn  vss 0.110f
C49 a2  vss 0.086f
C50 b   vss 0.081f
.ends
