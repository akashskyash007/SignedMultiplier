* Spice description of a2_x2
* Spice driver version 134999461
* Date  5/01/2008 at 14:59:11
* ssxlib 0.13um values
.subckt a2_x2 i0 i1 q vdd vss
Mtr_00001 sig2  i0    sig3  vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 vss   sig2  q     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00003 sig3  i1    vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00004 q     sig2  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00005 vdd   i1    sig2  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00006 sig2  i0    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C5  i0    vss   0.584f
C4  i1    vss   1.120f
C6  q     vss   0.815f
C2  sig2  vss   0.926f
.ends
