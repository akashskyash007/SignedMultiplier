.subckt oai21_x2 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from oai21_x2.ext -        technology: scmos
m00 vdd b  z   vdd p w=2.09u l=0.13u ad=0.707117p pd=3.46333u as=0.5962p   ps=3.42667u
m01 w1  a1 vdd vdd p w=2.09u l=0.13u ad=0.32395p  pd=2.4u     as=0.707117p ps=3.46333u
m02 z   a2 w1  vdd p w=2.09u l=0.13u ad=0.5962p   pd=3.42667u as=0.32395p  ps=2.4u    
m03 w2  a2 z   vdd p w=2.09u l=0.13u ad=0.32395p  pd=2.4u     as=0.5962p   ps=3.42667u
m04 vdd a1 w2  vdd p w=2.09u l=0.13u ad=0.707117p pd=3.46333u as=0.32395p  ps=2.4u    
m05 n3  b  z   vss n w=1.76u l=0.13u ad=0.4664p   pd=2.46667u as=0.59345p  ps=4.38u   
m06 vss a1 n3  vss n w=1.76u l=0.13u ad=0.6358p   pd=3.655u   as=0.4664p   ps=2.46667u
m07 n3  a2 vss vss n w=0.88u l=0.13u ad=0.2332p   pd=1.23333u as=0.3179p   ps=1.8275u 
m08 vss a2 n3  vss n w=0.88u l=0.13u ad=0.3179p   pd=1.8275u  as=0.2332p   ps=1.23333u
C0  a2  vdd 0.020f
C1  b   n3  0.013f
C2  z   vdd 0.082f
C3  a1  n3  0.068f
C4  a2  w2  0.020f
C5  z   w1  0.013f
C6  a2  n3  0.007f
C7  vdd w1  0.010f
C8  z   n3  0.018f
C9  vdd w2  0.010f
C10 b   a1  0.150f
C11 b   a2  0.017f
C12 b   z   0.134f
C13 a1  a2  0.254f
C14 a1  z   0.008f
C15 b   vdd 0.033f
C16 b   w1  0.010f
C17 a2  z   0.078f
C18 a1  vdd 0.037f
C19 n3  vss 0.124f
C20 w2  vss 0.013f
C21 w1  vss 0.012f
C23 z   vss 0.124f
C24 a2  vss 0.172f
C25 a1  vss 0.222f
C26 b   vss 0.127f
.ends
