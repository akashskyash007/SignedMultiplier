.subckt an4_x3 a b c d vdd vss z
*04-JAN-08 SPICE3       file   created      from an4_x3.ext -        technology: scmos
m00 z   zn vdd vdd p w=1.43u  l=0.13u ad=0.37895p  pd=1.96u    as=0.473985p ps=2.535u  
m01 vdd zn z   vdd p w=1.43u  l=0.13u ad=0.473985p pd=2.535u   as=0.37895p  ps=1.96u   
m02 zn  a  vdd vdd p w=1.595u l=0.13u ad=0.422675p pd=2.125u   as=0.528676p ps=2.8275u 
m03 vdd b  zn  vdd p w=1.595u l=0.13u ad=0.528676p pd=2.8275u  as=0.422675p ps=2.125u  
m04 zn  c  vdd vdd p w=1.595u l=0.13u ad=0.422675p pd=2.125u   as=0.528676p ps=2.8275u 
m05 vdd d  zn  vdd p w=1.595u l=0.13u ad=0.528676p pd=2.8275u  as=0.422675p ps=2.125u  
m06 vss zn z   vss n w=1.43u  l=0.13u ad=0.582907p pd=2.26068u as=0.506p    ps=3.72u   
m07 w1  a  vss vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.739843p ps=2.86932u
m08 w2  b  w1  vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.281325p ps=2.125u  
m09 w3  c  w2  vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.281325p ps=2.125u  
m10 zn  d  w3  vss n w=1.815u l=0.13u ad=0.608025p pd=4.49u    as=0.281325p ps=2.125u  
C0  w4 b   0.022f
C1  w5 c   0.010f
C2  w6 d   0.011f
C3  w7 vdd 0.034f
C4  zn a   0.244f
C5  w2 w5  0.002f
C6  w4 c   0.011f
C7  w5 d   0.002f
C8  w1 w5  0.002f
C9  zn b   0.110f
C10 z  vdd 0.053f
C11 w2 w4  0.006f
C12 w4 d   0.022f
C13 w1 w4  0.008f
C14 zn c   0.013f
C15 a  b   0.174f
C16 z  w7  0.016f
C17 w3 w4  0.006f
C18 w4 vdd 0.072f
C19 w2 zn  0.010f
C20 a  c   0.034f
C21 zn d   0.016f
C22 z  w6  0.009f
C23 w1 zn  0.010f
C24 w7 w4  0.166f
C25 w3 zn  0.010f
C26 zn vdd 0.221f
C27 b  c   0.226f
C28 z  w5  0.010f
C29 w6 w4  0.166f
C30 w7 zn  0.054f
C31 w2 b   0.016f
C32 a  vdd 0.021f
C33 b  d   0.003f
C34 z  w4  0.026f
C35 w1 b   0.009f
C36 w5 w4  0.166f
C37 w7 a   0.001f
C38 w6 zn  0.014f
C39 w3 b   0.010f
C40 b  vdd 0.010f
C41 c  d   0.151f
C42 z  zn  0.130f
C43 w7 b   0.001f
C44 w5 zn  0.021f
C45 w6 a   0.012f
C46 w3 c   0.004f
C47 c  vdd 0.010f
C48 w7 c   0.001f
C49 w4 zn  0.091f
C50 w5 a   0.002f
C51 d  vdd 0.032f
C52 w4 a   0.017f
C53 w5 b   0.009f
C54 w6 c   0.026f
C55 w7 d   0.002f
C56 w4 vss 0.954f
C57 w5 vss 0.175f
C58 w6 vss 0.172f
C59 w7 vss 0.149f
C60 w3 vss 0.010f
C61 w2 vss 0.010f
C62 w1 vss 0.010f
C63 z  vss 0.044f
C65 d  vss 0.099f
C66 c  vss 0.090f
C67 b  vss 0.076f
C68 a  vss 0.083f
C69 zn vss 0.336f
.ends
