.subckt nr3abv0x05 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from nr3abv0x05.ext -        technology: scmos
m00 w1  c  z   vdd p w=1.1u  l=0.13u ad=0.14025p  pd=1.355u   as=0.37015p  ps=2.95u   
m01 vdd nd w1  vdd p w=1.1u  l=0.13u ad=0.42075p  pd=3.02273u as=0.14025p  ps=1.355u  
m02 nd  a  vdd vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.25245p  ps=1.81364u
m03 vdd b  nd  vdd p w=0.66u l=0.13u ad=0.25245p  pd=1.81364u as=0.1386p   ps=1.08u   
m04 z   c  vss vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.14025p  ps=1.21364u
m05 vss nd z   vss n w=0.33u l=0.13u ad=0.14025p  pd=1.21364u as=0.0693p   ps=0.75u   
m06 w2  a  vss vss n w=0.55u l=0.13u ad=0.070125p pd=0.805u   as=0.23375p  ps=2.02273u
m07 nd  b  w2  vss n w=0.55u l=0.13u ad=0.18205p  pd=1.85u    as=0.070125p ps=0.805u  
C0  c   a   0.020f
C1  nd  a   0.170f
C2  z   a   0.004f
C3  nd  b   0.089f
C4  vdd c   0.032f
C5  a   b   0.089f
C6  vdd nd  0.007f
C7  vdd z   0.018f
C8  vdd w1  0.003f
C9  c   nd  0.160f
C10 c   z   0.114f
C11 nd  z   0.005f
C12 c   w1  0.008f
C13 vdd b   0.072f
C14 w2  vss 0.006f
C15 b   vss 0.111f
C16 a   vss 0.125f
C17 w1  vss 0.006f
C18 z   vss 0.275f
C19 nd  vss 0.172f
C20 c   vss 0.110f
.ends
