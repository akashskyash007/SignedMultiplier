.subckt vsstie vdd vss z
*10-JAN-08 SPICE3       file   created      from vsstie.ext -        technology: scmos
m00 w1  z  vdd vdd p w=1.43u l=0.13u ad=0.37895p pd=1.96u as=0.53625p ps=3.61u
m01 vdd z  w1  vdd p w=1.43u l=0.13u ad=0.53625p pd=3.61u as=0.37895p ps=1.96u
m02 z   w1 vss vss n w=0.99u l=0.13u ad=0.26235p pd=1.52u as=0.37125p ps=2.73u
m03 vss w1 z   vss n w=0.99u l=0.13u ad=0.37125p pd=2.73u as=0.26235p ps=1.52u
C0 vdd z   0.093f
C1 vdd w1  0.061f
C2 z   w1  0.267f
C3 w1  vss 0.288f
C4 z   vss 0.369f
.ends
