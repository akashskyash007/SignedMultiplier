.subckt aoi21a2bv0x05 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from aoi21a2bv0x05.ext -        technology: scmos
m00 vdd a2  a2n vdd p w=0.66u  l=0.13u ad=0.235832p  pd=1.515u    as=0.2112p    ps=2.07u    
m01 bn  b   vdd vdd p w=0.66u  l=0.13u ad=0.2112p    pd=2.07u     as=0.235832p  ps=1.515u   
m02 n1  bn  z   vdd p w=0.88u  l=0.13u ad=0.22715p   pd=1.70333u  as=0.2695p    ps=2.51u    
m03 vdd a2n n1  vdd p w=0.88u  l=0.13u ad=0.314443p  pd=2.02u     as=0.22715p   ps=1.70333u 
m04 n1  a1  vdd vdd p w=0.88u  l=0.13u ad=0.22715p   pd=1.70333u  as=0.314443p  ps=2.02u    
m05 bn  b   vss vss n w=0.33u  l=0.13u ad=0.12375p   pd=1.41u     as=0.275484p  ps=2.0664u  
m06 z   bn  vss vss n w=0.33u  l=0.13u ad=0.0706962p pd=0.743077u as=0.275484p  ps=2.0664u  
m07 vss a2  a2n vss n w=0.33u  l=0.13u ad=0.275484p  pd=2.0664u   as=0.12375p   ps=1.41u    
m08 w1  a2n z   vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u     as=0.0824789p ps=0.866923u
m09 vss a1  w1  vss n w=0.385u l=0.13u ad=0.321398p  pd=2.4108u   as=0.0490875p ps=0.64u    
C0  a1  z   0.007f
C1  a2n bn  0.082f
C2  a2n z   0.083f
C3  a1  n1  0.052f
C4  vdd a2  0.066f
C5  bn  z   0.116f
C6  a2n n1  0.006f
C7  vdd b   0.003f
C8  a2n w1  0.012f
C9  vdd a1  0.009f
C10 z   n1  0.036f
C11 vdd a2n 0.007f
C12 a2  b   0.115f
C13 vdd bn  0.005f
C14 a2  a2n 0.066f
C15 a2  bn  0.023f
C16 b   a2n 0.069f
C17 vdd n1  0.043f
C18 b   bn  0.084f
C19 a1  a2n 0.077f
C20 b   z   0.008f
C21 n1  vss 0.049f
C22 z   vss 0.059f
C23 bn  vss 0.123f
C24 a2n vss 0.559f
C25 a1  vss 0.106f
C26 b   vss 0.122f
C27 a2  vss 0.099f
.ends
