* Spice description of no3_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:18:51
* sxlib 0.13um values
.subckt no3_x1 i0 i1 i2 nq vdd vss
Mtr_00001 vss   i0    nq    vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 nq    i2    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 nq    i1    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00004 vdd   i2    sig5  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00005 sig3  i1    nq    vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00006 sig5  i0    sig3  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C7  i0    vss   0.932f
C6  i1    vss   0.915f
C8  i2    vss   1.050f
C1  nq    vss   0.988f
.ends
