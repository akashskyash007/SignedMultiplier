* Spice description of nd2ab_x2
* Spice driver version 134999461
* Date  4/01/2008 at 19:02:09
* vxlib 0.13um values
.subckt nd2ab_x2 a b vdd vss z
M1a sig5  a     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M1b vdd   b     bn    vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M1z vdd   sig5  z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2a vss   a     sig5  vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M2b bn    b     vss   vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M2z z     bn    vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3z n1    sig5  vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M4z z     bn    n1    vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C8  a     vss   0.813f
C3  bn    vss   0.958f
C7  b     vss   0.713f
C5  sig5  vss   0.760f
C1  z     vss   0.737f
.ends
