.subckt vddtie vdd vss z
*01-JAN-08 SPICE3       file   created      from vddtie.ext -        technology: scmos
m00 z vss vdd vdd p w=1.045u l=0.13u ad=0.44935p pd=2.95u as=0.73975p ps=4.27u
m01 z vss vss vss n w=0.55u  l=0.13u ad=0.2365p  pd=1.96u as=0.52085p ps=3.39u
C0 vdd z   0.064f
C1 z   vss 0.201f
.ends
