* Spice description of iv1v0x4
* Spice driver version 134999461
* Date 10/01/2008 at 14:50:26
* rgalib 0.13um values
.subckt iv1v0x4 a vdd vss z
Mtr_00001 vss   a     z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 z     a     vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 vdd   a     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00004 z     a     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
C3  a     vss   1.161f
C1  z     vss   1.449f
.ends
