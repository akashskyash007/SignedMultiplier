* Spice description of nd2v5x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:51:51
* vsclib 0.13um values
.subckt nd2v5x2 a b vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 vss   a     sig3  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M03 z     b     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 sig3  b     z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
C4  a     vss   0.597f
C5  b     vss   0.333f
C1  z     vss   0.594f
.ends
