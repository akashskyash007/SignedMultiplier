.subckt nd2v5x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v5x2.ext -        technology: scmos
m00 z   b vdd vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u  as=0.61985p  ps=3.885u
m01 vdd a z   vdd p w=1.54u l=0.13u ad=0.61985p  pd=3.885u as=0.3234p   ps=1.96u 
m02 w1  b z   vss n w=0.99u l=0.13u ad=0.126225p pd=1.245u as=0.29865p  ps=2.73u 
m03 vss a w1  vss n w=0.99u l=0.13u ad=0.48015p  pd=2.95u  as=0.126225p ps=1.245u
C0  b   a   0.137f
C1  b   vdd 0.007f
C2  b   z   0.078f
C3  a   vdd 0.027f
C4  b   w1  0.007f
C5  a   z   0.004f
C6  vdd z   0.091f
C7  w1  vss 0.008f
C8  z   vss 0.214f
C10 a   vss 0.110f
C11 b   vss 0.083f
.ends
