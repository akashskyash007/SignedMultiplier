.subckt bf1v0x8 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v0x8.ext -        technology: scmos
m00 z   an vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.85u    as=0.378415p ps=2.4302u  
m01 vdd an z   vdd p w=1.43u  l=0.13u ad=0.378415p pd=2.4302u  as=0.3003p   ps=1.85u    
m02 z   an vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.85u    as=0.378415p ps=2.4302u  
m03 vdd an z   vdd p w=1.43u  l=0.13u ad=0.378415p pd=2.4302u  as=0.3003p   ps=1.85u    
m04 an  a  vdd vdd p w=1.43u  l=0.13u ad=0.316762p pd=2.23721u as=0.378415p ps=2.4302u  
m05 vdd a  an  vdd p w=0.935u l=0.13u ad=0.247425p pd=1.58898u as=0.207113p ps=1.46279u 
m06 z   an vss vss n w=0.715u l=0.13u ad=0.15015p  pd=1.135u   as=0.191572p ps=1.50453u 
m07 vss an z   vss n w=0.715u l=0.13u ad=0.191572p pd=1.50453u as=0.15015p  ps=1.135u   
m08 z   an vss vss n w=0.715u l=0.13u ad=0.15015p  pd=1.135u   as=0.191572p ps=1.50453u 
m09 vss an z   vss n w=0.715u l=0.13u ad=0.191572p pd=1.50453u as=0.15015p  ps=1.135u   
m10 an  a  vss vss n w=0.715u l=0.13u ad=0.155279p pd=1.28304u as=0.191572p ps=1.50453u 
m11 vss a  an  vss n w=0.55u  l=0.13u ad=0.147363p pd=1.15733u as=0.119446p ps=0.986957u
C0 vdd z   0.031f
C1 an  a   0.149f
C2 an  z   0.178f
C3 vdd an  0.034f
C4 vdd a   0.027f
C5 z   vss 0.299f
C6 a   vss 0.164f
C7 an  vss 0.350f
.ends
