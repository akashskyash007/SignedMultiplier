.subckt noa22_x1 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa22_x1.ext -        technology: scmos
m00 nq  i0 w1  vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u    as=0.69715p ps=3.55667u
m01 w1  i1 nq  vdd p w=2.19u l=0.13u ad=0.69715p pd=3.55667u as=0.58035p ps=2.72u   
m02 vdd i2 w1  vdd p w=2.19u l=0.13u ad=0.93075p pd=5.23u    as=0.69715p ps=3.55667u
m03 w2  i0 vss vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u    as=0.46325p ps=3.03u   
m04 nq  i1 w2  vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u    as=0.28885p ps=1.62u   
m05 vss i2 nq  vss n w=1.09u l=0.13u ad=0.46325p pd=3.03u    as=0.28885p ps=1.62u   
C0  vdd w1  0.099f
C1  i0  i1  0.221f
C2  vdd nq  0.019f
C3  i0  w1  0.014f
C4  i1  i2  0.096f
C5  i1  w1  0.005f
C6  i1  nq  0.146f
C7  i2  w1  0.010f
C8  i1  w2  0.015f
C9  i2  nq  0.140f
C10 w1  nq  0.095f
C11 vdd i0  0.010f
C12 vdd i1  0.010f
C13 vdd i2  0.113f
C14 w2  vss 0.027f
C15 nq  vss 0.128f
C16 w1  vss 0.076f
C17 i2  vss 0.210f
C18 i1  vss 0.154f
C19 i0  vss 0.158f
.ends
