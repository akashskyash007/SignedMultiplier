.subckt nd2v0x05 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v0x05.ext -        technology: scmos
m00 z   b vdd vdd p w=0.44u  l=0.13u ad=0.0924p    pd=0.86u  as=0.397925p  ps=3.005u
m01 vdd a z   vdd p w=0.44u  l=0.13u ad=0.397925p  pd=3.005u as=0.0924p    ps=0.86u 
m02 w1  b z   vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u  as=0.144375p  ps=1.52u 
m03 vss a w1  vss n w=0.385u l=0.13u ad=0.33495p   pd=2.51u  as=0.0490875p ps=0.64u 
C0 b   a   0.066f
C1 b   z   0.032f
C2 a   z   0.004f
C3 vdd b   0.076f
C4 vdd a   0.010f
C5 vdd z   0.014f
C6 w1  vss 0.001f
C7 z   vss 0.082f
C8 a   vss 0.109f
C9 b   vss 0.117f
.ends
