* Spice description of iv1_x2
* Spice driver version 134999461
* Date  4/01/2008 at 19:00:01
* vsxlib 0.13um values
.subckt iv1_x2 a vdd vss z
M1  vdd   a     z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2  z     a     vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C3  a     vss   0.591f
C1  z     vss   0.694f
.ends
