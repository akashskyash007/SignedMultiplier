.subckt xaoi21v0x1 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from xaoi21v0x1.ext -        technology: scmos
m00 bn  b  vdd vdd p w=1.54u  l=0.13u ad=0.4444p   pd=3.83u    as=0.53515p  ps=3.005u  
m01 z   b  an  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.363733p ps=2.58333u
m02 w1  an z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m03 vdd bn w1  vdd p w=1.54u  l=0.13u ad=0.53515p  pd=3.005u   as=0.19635p  ps=1.795u  
m04 an  a2 vdd vdd p w=1.54u  l=0.13u ad=0.363733p pd=2.58333u as=0.53515p  ps=3.005u  
m05 vdd a1 an  vdd p w=1.54u  l=0.13u ad=0.53515p  pd=3.005u   as=0.363733p ps=2.58333u
m06 bn  b  vss vss n w=0.715u l=0.13u ad=0.15015p  pd=1.135u   as=0.268125p ps=2.08u   
m07 z   an bn  vss n w=0.715u l=0.13u ad=0.236665p pd=2.17533u as=0.15015p  ps=1.135u  
m08 an  bn z   vss n w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.309485p ps=2.84467u
m09 w2  a2 an  vss n w=0.935u l=0.13u ad=0.119213p pd=1.19u    as=0.19635p  ps=1.355u  
m10 vss a1 w2  vss n w=0.935u l=0.13u ad=0.350625p pd=2.72u    as=0.119213p ps=1.19u   
C0  an  a1  0.016f
C1  b   vdd 0.028f
C2  bn  a2  0.084f
C3  b   z   0.013f
C4  an  vdd 0.188f
C5  an  z   0.121f
C6  bn  vdd 0.012f
C7  a2  a1  0.155f
C8  bn  z   0.163f
C9  an  w1  0.008f
C10 a2  vdd 0.027f
C11 bn  w1  0.014f
C12 a1  vdd 0.007f
C13 vdd z   0.007f
C14 b   an  0.097f
C15 a1  w2  0.009f
C16 vdd w1  0.004f
C17 b   bn  0.050f
C18 an  bn  0.323f
C19 an  a2  0.114f
C20 w2  vss 0.009f
C21 w1  vss 0.006f
C22 z   vss 0.143f
C24 a1  vss 0.134f
C25 a2  vss 0.095f
C26 bn  vss 0.187f
C27 an  vss 0.223f
C28 b   vss 0.202f
.ends
