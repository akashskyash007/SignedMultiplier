.subckt nd2_x2 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nd2_x2.ext -        technology: scmos
m00 z   b vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=1.04033p  ps=5.26u 
m01 vdd a z   vdd p w=2.145u l=0.13u ad=1.04033p  pd=5.26u  as=0.568425p ps=2.675u
m02 w1  b z   vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u as=0.608025p ps=4.49u 
m03 vss a w1  vss n w=1.815u l=0.13u ad=0.880275p pd=4.6u   as=0.281325p ps=2.125u
C0  b   a   0.209f
C1  b   vdd 0.020f
C2  b   z   0.108f
C3  a   vdd 0.010f
C4  a   z   0.012f
C5  a   w1  0.004f
C6  vdd z   0.110f
C7  w1  vss 0.020f
C8  z   vss 0.139f
C10 a   vss 0.146f
C11 b   vss 0.110f
.ends
