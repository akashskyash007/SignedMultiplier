.subckt oa2a22_x2 i0 i1 i2 i3 q vdd vss
*05-JAN-08 SPICE3       file   created      from oa2a22_x2.ext -        technology: scmos
m00 w1  i0 w2  vdd p w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.37605p  ps=2.325u  
m01 w2  i1 w1  vdd p w=1.09u l=0.13u ad=0.37605p  pd=2.325u   as=0.28885p  ps=1.62u   
m02 vdd i2 w2  vdd p w=1.09u l=0.13u ad=0.411369p pd=2.33215u as=0.37605p  ps=2.325u  
m03 w2  i3 vdd vdd p w=1.09u l=0.13u ad=0.37605p  pd=2.325u   as=0.411369p ps=2.33215u
m04 q   w1 vdd vdd p w=2.19u l=0.13u ad=0.93075p  pd=5.23u    as=0.826512p ps=4.6857u 
m05 w3  i0 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.299576p ps=2.15253u
m06 w1  i1 w3  vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.1431p   ps=1.07u   
m07 w4  i2 w1  vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.1431p   ps=1.07u   
m08 vss i3 w4  vss n w=0.54u l=0.13u ad=0.299576p pd=2.15253u as=0.1431p   ps=1.07u   
m09 q   w1 vss vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.604699p ps=4.34493u
C0  w1  i2  0.113f
C1  vdd w2  0.140f
C2  i0  i1  0.201f
C3  i1  w3  0.015f
C4  w1  i3  0.014f
C5  w1  w2  0.124f
C6  i1  i2  0.076f
C7  i2  w4  0.015f
C8  i0  w2  0.005f
C9  i1  w2  0.005f
C10 i2  i3  0.201f
C11 i2  w2  0.005f
C12 vdd w1  0.061f
C13 vdd q   0.033f
C14 i3  w2  0.005f
C15 vdd i0  0.002f
C16 vdd i1  0.002f
C17 w1  q   0.075f
C18 vdd i2  0.002f
C19 w1  i1  0.114f
C20 vdd i3  0.002f
C21 w4  vss 0.006f
C22 w3  vss 0.006f
C23 q   vss 0.122f
C24 w2  vss 0.066f
C25 i3  vss 0.167f
C26 i2  vss 0.167f
C27 i1  vss 0.167f
C28 i0  vss 0.168f
C29 w1  vss 0.213f
.ends
