.subckt nd2v5x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v5x1.ext -        technology: scmos
m00 z   b vdd vdd p w=1.045u l=0.13u ad=0.21945p pd=1.465u as=0.4675p  ps=3.06u 
m01 vdd a z   vdd p w=1.045u l=0.13u ad=0.4675p  pd=3.06u  as=0.21945p ps=1.465u
m02 w1  b z   vss n w=0.66u  l=0.13u ad=0.08415p pd=0.915u as=0.2112p  ps=2.07u 
m03 vss a w1  vss n w=0.66u  l=0.13u ad=0.429p   pd=2.62u  as=0.08415p ps=0.915u
C0 b   a   0.119f
C1 b   z   0.079f
C2 a   z   0.008f
C3 vdd b   0.003f
C4 vdd z   0.087f
C5 w1  vss 0.008f
C6 z   vss 0.184f
C7 a   vss 0.135f
C8 b   vss 0.101f
.ends
