* Spice description of one_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:36:37
* sxlib 0.13um values
.subckt one_x0 q vdd vss
Mtr_00001 q     vss   vdd   vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
C1  q     vss   0.731f
.ends
