* Spice description of vfeed6
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:46
* vxlib 0.13um values
.subckt vfeed6 vdd vss
.ends
