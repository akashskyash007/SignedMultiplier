.subckt bf1v0x1 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v0x1.ext -        technology: scmos
m00 vdd an z   vdd p w=0.99u  l=0.13u ad=0.4257p   pd=2.59548u as=0.341p    ps=2.73u    
m01 an  a  vdd vdd p w=0.715u l=0.13u ad=0.225775p pd=2.18u    as=0.30745p  ps=1.87452u 
m02 vss an z   vss n w=0.495u l=0.13u ad=0.135979p pd=1.08529u as=0.167475p ps=1.74u    
m03 an  a  vss vss n w=0.44u  l=0.13u ad=0.1529p   pd=1.63u    as=0.120871p ps=0.964706u
C0 z   a   0.023f
C1 vdd z   0.009f
C2 vdd a   0.052f
C3 an  z   0.026f
C4 an  a   0.066f
C5 a   vss 0.087f
C6 z   vss 0.134f
C7 an  vss 0.125f
.ends
