* Spice description of aon21_x1
* Spice driver version 134999461
* Date  4/01/2008 at 18:51:54
* vxlib 0.13um values
.subckt aon21_x1 a1 a2 b vdd vss z
M1  vdd   a1    sig5  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M2  sig5  a2    vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M3_1 z     zn    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M3  zn    b     sig5  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M4  vss   a1    n1    vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M5_2 vss   zn    z     vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M5  n1    a2    zn    vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M6  zn    b     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C8  a1    vss   0.880f
C7  a2    vss   0.769f
C9  b     vss   0.839f
C5  sig5  vss   0.184f
C1  zn    vss   0.890f
C4  z     vss   0.591f
.ends
