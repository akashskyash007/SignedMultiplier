.subckt oan21_x2 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from oan21_x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=2.09u  l=0.13u ad=0.755013p pd=4.06917u as=0.6809p   ps=5.04u   
m01 zn  b  vdd vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.8069u  as=0.397375p ps=2.14167u
m02 w1  a2 zn  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.55385p  ps=3.4331u 
m03 vdd a1 w1  vdd p w=2.09u  l=0.13u ad=0.755013p pd=4.06917u as=0.32395p  ps=2.4u    
m04 z   zn vss vss n w=1.045u l=0.13u ad=0.403975p pd=2.95u    as=0.371271p ps=2.62057u
m05 n2  b  zn  vss n w=0.935u l=0.13u ad=0.290125p pd=1.88667u as=0.374825p ps=2.73u   
m06 vss a2 n2  vss n w=0.935u l=0.13u ad=0.33219p  pd=2.34472u as=0.290125p ps=1.88667u
m07 n2  a1 vss vss n w=0.935u l=0.13u ad=0.290125p pd=1.88667u as=0.33219p  ps=2.34472u
C0  zn  w2  0.006f
C1  a2  n2  0.010f
C2  a1  w1  0.012f
C3  w3  zn  0.042f
C4  w4  w3  0.166f
C5  zn  w5  0.023f
C6  a2  w2  0.002f
C7  a1  n2  0.007f
C8  w3  a2  0.013f
C9  vdd zn  0.050f
C10 a2  w5  0.011f
C11 a1  w2  0.002f
C12 w3  a1  0.018f
C13 vdd a2  0.010f
C14 a1  w5  0.011f
C15 z   w2  0.004f
C16 b   n2  0.073f
C17 w3  z   0.023f
C18 vdd a1  0.065f
C19 w4  zn  0.020f
C20 z   w5  0.030f
C21 b   w2  0.001f
C22 w3  b   0.018f
C23 zn  a2  0.013f
C24 vdd z   0.015f
C25 w4  a2  0.029f
C26 b   w5  0.001f
C27 w1  w2  0.005f
C28 w3  w1  0.008f
C29 zn  a1  0.016f
C30 w1  w5  0.001f
C31 w3  n2  0.040f
C32 zn  z   0.145f
C33 vdd w1  0.009f
C34 a2  a1  0.224f
C35 w4  z   0.009f
C36 w3  w2  0.166f
C37 zn  b   0.151f
C38 w4  b   0.011f
C39 w3  w5  0.166f
C40 vdd w2  0.024f
C41 a2  b   0.141f
C42 w3  vdd 0.054f
C43 vdd w5  0.008f
C44 zn  n2  0.007f
C45 a2  w1  0.017f
C46 a1  b   0.002f
C47 w3  vss 0.990f
C48 w4  vss 0.172f
C49 w5  vss 0.163f
C50 w2  vss 0.172f
C51 n2  vss 0.086f
C52 b   vss 0.093f
C53 z   vss 0.059f
C54 a1  vss 0.068f
C55 a2  vss 0.087f
C56 zn  vss 0.109f
.ends
