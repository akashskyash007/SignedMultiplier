.subckt nd2v0x2 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from nd2v0x2.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 vdd b z   vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 w1  a vss vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m03 z   b w1  vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0  a   z   0.091f
C1  a   b   0.089f
C2  z   b   0.126f
C3  z   w1  0.022f
C4  vdd a   0.038f
C5  vdd z   0.018f
C6  vdd b   0.038f
C7  w1  vss 0.023f
C8  b   vss 0.153f
C9  z   vss 0.084f
C10 a   vss 0.178f
.ends
