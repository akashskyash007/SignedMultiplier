.subckt nr2_x2 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2_x2.ext -        technology: scmos
m00 w1  a vdd vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=1.04033p  ps=5.26u 
m01 z   b w1  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.332475p ps=2.455u
m02 w2  b z   vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=0.568425p ps=2.675u
m03 vdd a w2  vdd p w=2.145u l=0.13u ad=1.04033p  pd=5.26u  as=0.332475p ps=2.455u
m04 z   a vss vss n w=1.155u l=0.13u ad=0.306075p pd=1.685u as=0.560175p ps=3.28u 
m05 vss b z   vss n w=1.155u l=0.13u ad=0.560175p pd=3.28u  as=0.306075p ps=1.685u
C0  a   b   0.303f
C1  a   vdd 0.020f
C2  b   vdd 0.020f
C3  a   z   0.099f
C4  b   z   0.042f
C5  vdd w1  0.010f
C6  b   w2  0.017f
C7  vdd z   0.053f
C8  w1  z   0.012f
C9  vdd w2  0.010f
C10 w2  vss 0.012f
C11 z   vss 0.234f
C12 w1  vss 0.012f
C14 b   vss 0.136f
C15 a   vss 0.200f
.ends
