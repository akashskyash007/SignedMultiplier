.subckt nr2av0x3 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2av0x3.ext -        technology: scmos
m00 w1  b  z   vdd p w=1.375u l=0.13u ad=0.175313p pd=1.63u    as=0.340175p ps=2.36333u
m01 vdd an w1  vdd p w=1.375u l=0.13u ad=0.309308p pd=1.84951u as=0.175313p ps=1.63u   
m02 w2  an vdd vdd p w=1.375u l=0.13u ad=0.175313p pd=1.63u    as=0.309308p ps=1.84951u
m03 z   b  w2  vdd p w=1.375u l=0.13u ad=0.340175p pd=2.36333u as=0.175313p ps=1.63u   
m04 w3  b  z   vdd p w=1.375u l=0.13u ad=0.175313p pd=1.63u    as=0.340175p ps=2.36333u
m05 vdd an w3  vdd p w=1.375u l=0.13u ad=0.309308p pd=1.84951u as=0.175313p ps=1.63u   
m06 an  a  vdd vdd p w=1.54u  l=0.13u ad=0.48675p  pd=3.83u    as=0.346425p ps=2.07146u
m07 z   b  vss vss n w=1.1u   l=0.13u ad=0.231p    pd=1.52u    as=0.525657p ps=3.44074u
m08 vss an z   vss n w=1.1u   l=0.13u ad=0.525657p pd=3.44074u as=0.231p    ps=1.52u   
m09 an  a  vss vss n w=0.77u  l=0.13u ad=0.28875p  pd=2.29u    as=0.36796p  ps=2.40852u
C0  vdd w2  0.004f
C1  b   an  0.345f
C2  vdd w3  0.004f
C3  b   a   0.028f
C4  b   z   0.183f
C5  an  a   0.166f
C6  an  z   0.046f
C7  b   vdd 0.021f
C8  an  vdd 0.026f
C9  z   w1  0.009f
C10 a   vdd 0.009f
C11 z   vdd 0.101f
C12 a   w3  0.002f
C13 z   w2  0.009f
C14 w1  vdd 0.004f
C15 w3  vss 0.010f
C16 w2  vss 0.007f
C18 w1  vss 0.008f
C19 z   vss 0.141f
C20 a   vss 0.099f
C21 an  vss 0.302f
C22 b   vss 0.469f
.ends
