.subckt nr2av0x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2av0x2.ext -        technology: scmos
m00 w1  an vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.45045p  ps=2.751u  
m01 z   b  w1  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.19635p  ps=1.795u  
m02 w2  b  z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m03 vdd an w2  vdd p w=1.54u  l=0.13u ad=0.45045p  pd=2.751u   as=0.19635p  ps=1.795u  
m04 an  a  vdd vdd p w=1.32u  l=0.13u ad=0.42845p  pd=3.39u    as=0.3861p   ps=2.358u  
m05 z   an vss vss n w=0.825u l=0.13u ad=0.17325p  pd=1.245u   as=0.405527p ps=2.53214u
m06 vss b  z   vss n w=0.825u l=0.13u ad=0.405527p pd=2.53214u as=0.17325p  ps=1.245u  
m07 an  a  vss vss n w=0.66u  l=0.13u ad=0.2112p   pd=2.07u    as=0.324421p ps=2.02571u
C0  an  z   0.133f
C1  b   w1  0.006f
C2  b   z   0.127f
C3  vdd w1  0.004f
C4  vdd z   0.021f
C5  an  a   0.147f
C6  vdd w2  0.004f
C7  b   a   0.007f
C8  vdd a   0.005f
C9  z   w2  0.009f
C10 an  b   0.224f
C11 an  vdd 0.020f
C12 b   vdd 0.017f
C13 a   vss 0.133f
C14 w2  vss 0.008f
C15 z   vss 0.085f
C16 w1  vss 0.009f
C18 b   vss 0.099f
C19 an  vss 0.436f
.ends
