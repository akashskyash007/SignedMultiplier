.subckt vfeed8 vdd vss
*01-JAN-08 SPICE3       file   created      from vfeed8.ext -        technology: scmos
.ends
