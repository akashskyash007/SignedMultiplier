.subckt no2_x4 i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from no2_x4.ext -        technology: scmos
m00 w1  i1 w2  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.8987p   ps=5.04u   
m01 vdd i0 w1  vdd p w=2.09u  l=0.13u ad=0.663729p pd=3.05118u as=0.32395p  ps=2.4u    
m02 nq  w3 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.681195p ps=3.13147u
m03 vdd w3 nq  vdd p w=2.145u l=0.13u ad=0.681195p pd=3.13147u as=0.568425p ps=2.675u  
m04 w3  w2 vdd vdd p w=1.1u   l=0.13u ad=0.473p    pd=3.06u    as=0.349331p ps=1.60588u
m05 w2  i1 vss vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.200912p ps=1.40882u
m06 vss i0 w2  vss n w=0.55u  l=0.13u ad=0.200912p pd=1.40882u as=0.14575p  ps=1.08u   
m07 nq  w3 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.381732p ps=2.67676u
m08 vss w3 nq  vss n w=1.045u l=0.13u ad=0.381732p pd=2.67676u as=0.276925p ps=1.575u  
m09 w3  w2 vss vss n w=0.55u  l=0.13u ad=0.2365p   pd=1.96u    as=0.200912p ps=1.40882u
C0  i0  w1  0.012f
C1  w3  w2  0.193f
C2  w3  nq  0.032f
C3  w2  w1  0.010f
C4  w2  nq  0.213f
C5  vdd i1  0.010f
C6  vdd i0  0.022f
C7  vdd w3  0.020f
C8  vdd w2  0.266f
C9  i1  i0  0.249f
C10 vdd w1  0.010f
C11 i1  w2  0.039f
C12 vdd nq  0.017f
C13 i0  w3  0.078f
C14 i0  w2  0.157f
C15 nq  vss 0.121f
C16 w1  vss 0.010f
C17 w2  vss 0.344f
C18 w3  vss 0.305f
C19 i0  vss 0.130f
C20 i1  vss 0.132f
.ends
