* Spice description of nd2v0x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:49:59
* wsclib 0.13um values
.subckt nd2v0x2 a b vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M02 vss   a     sig3  vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M03 z     b     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M04 sig3  b     z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C5  a     vss   0.560f
C4  b     vss   0.374f
C2  z     vss   0.594f
.ends
