.subckt mx2_x2 cmd i0 i1 q vdd vss
*05-JAN-08 SPICE3       file   created      from mx2_x2.ext -        technology: scmos
m00 vdd cmd w1  vdd p w=1.09u l=0.13u ad=0.49615p  pd=2.08418u as=0.46325p  ps=3.03u   
m01 w2  i0  vdd vdd p w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.49615p  ps=2.08418u
m02 w3  cmd w2  vdd p w=1.09u l=0.13u ad=0.40875p  pd=1.84u    as=0.16895p  ps=1.4u    
m03 w4  w1  w3  vdd p w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.40875p  ps=1.84u   
m04 vdd i1  w4  vdd p w=1.09u l=0.13u ad=0.49615p  pd=2.08418u as=0.16895p  ps=1.4u    
m05 q   w3  vdd vdd p w=2.19u l=0.13u ad=0.93075p  pd=5.23u    as=0.996851p ps=4.18747u
m06 vss cmd w1  vss n w=0.54u l=0.13u ad=0.256201p pd=1.24738u as=0.4055p   ps=3.03u   
m07 w5  i0  vss vss n w=0.54u l=0.13u ad=0.0837p   pd=0.85u    as=0.256201p ps=1.24738u
m08 w3  w1  w5  vss n w=0.54u l=0.13u ad=0.41535p  pd=2.28u    as=0.0837p   ps=0.85u   
m09 w6  cmd w3  vss n w=0.54u l=0.13u ad=0.0837p   pd=0.85u    as=0.41535p  ps=2.28u   
m10 vss i1  w6  vss n w=0.54u l=0.13u ad=0.256201p pd=1.24738u as=0.0837p   ps=0.85u   
m11 q   w3  vss vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.517147p ps=2.51786u
C0  w1  i1  0.136f
C1  vdd w3  0.021f
C2  vdd cmd 0.015f
C3  vdd i0  0.046f
C4  vdd w1  0.012f
C5  w3  cmd 0.181f
C6  vdd i1  0.108f
C7  w3  w1  0.101f
C8  cmd i0  0.296f
C9  cmd w1  0.046f
C10 w3  i1  0.024f
C11 vdd q   0.093f
C12 cmd i1  0.052f
C13 i0  w1  0.134f
C14 cmd w2  0.020f
C15 w6  vss 0.012f
C16 w5  vss 0.012f
C17 q   vss 0.133f
C18 w4  vss 0.010f
C19 w2  vss 0.006f
C20 i1  vss 0.194f
C21 w1  vss 0.439f
C22 i0  vss 0.152f
C23 cmd vss 0.339f
C24 w3  vss 0.228f
.ends
