* Spice description of vfeed6
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:58
* vsclib 0.13um values
.subckt vfeed6 vdd vss
.ends
