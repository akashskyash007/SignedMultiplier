.subckt nd2v3x3 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v3x3.ext -        technology: scmos
m00 z   b vdd vdd p w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.286344p ps=2.015u  
m01 vdd a z   vdd p w=0.935u l=0.13u ad=0.286344p pd=2.015u   as=0.19635p  ps=1.355u  
m02 z   a vdd vdd p w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.286344p ps=2.015u  
m03 vdd b z   vdd p w=0.935u l=0.13u ad=0.286344p pd=2.015u   as=0.19635p  ps=1.355u  
m04 w1  b z   vss n w=0.935u l=0.13u ad=0.119213p pd=1.19u    as=0.235144p ps=1.68807u
m05 vss a w1  vss n w=0.935u l=0.13u ad=0.291982p pd=1.85211u as=0.119213p ps=1.19u   
m06 w2  a vss vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.343509p ps=2.17895u
m07 z   b w2  vss n w=1.1u   l=0.13u ad=0.27664p  pd=1.98597u as=0.14025p  ps=1.355u  
m08 w3  b z   vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.27664p  ps=1.98597u
m09 vss a w3  vss n w=1.1u   l=0.13u ad=0.343509p pd=2.17895u as=0.14025p  ps=1.355u  
C0  b   w2  0.006f
C1  z   w1  0.009f
C2  z   w2  0.009f
C3  vdd b   0.008f
C4  vdd a   0.018f
C5  vdd z   0.134f
C6  b   a   0.447f
C7  b   z   0.230f
C8  a   z   0.077f
C9  w3  vss 0.012f
C10 w2  vss 0.009f
C11 w1  vss 0.005f
C12 z   vss 0.387f
C13 a   vss 0.250f
C14 b   vss 0.248f
.ends
