* Spice description of noa3ao322_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:25:03
* sxlib 0.13um values
.subckt noa3ao322_x1 i0 i1 i2 i3 i4 i5 i6 nq vdd vss
Mtr_00001 vss   i5    sig3  vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00002 sig3  i4    vss   vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00003 vss   i3    sig3  vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00004 sig3  i6    nq    vss n  L=0.12U  W=0.98U  AS=0.2597P   AD=0.2597P   PS=2.49U   PD=2.49U
Mtr_00005 nq    i2    sig4  vss n  L=0.12U  W=1.31U  AS=0.34715P  AD=0.34715P  PS=3.15U   PD=3.15U
Mtr_00006 sig4  i1    sig5  vss n  L=0.12U  W=1.31U  AS=0.34715P  AD=0.34715P  PS=3.15U   PD=3.15U
Mtr_00007 sig5  i0    vss   vss n  L=0.12U  W=1.31U  AS=0.34715P  AD=0.34715P  PS=3.15U   PD=3.15U
Mtr_00008 sig7  i0    vdd   vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00009 vdd   i1    sig7  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00010 sig7  i2    vdd   vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00011 sig7  i5    sig14 vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00012 sig14 i4    sig8  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00013 nq    i6    sig7  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00014 sig8  i3    nq    vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C11 i0    vss   0.766f
C10 i1    vss   0.800f
C12 i2    vss   0.699f
C13 i3    vss   0.565f
C16 i4    vss   0.699f
C15 i5    vss   0.665f
C9  i6    vss   0.654f
C2  nq    vss   0.764f
C3  sig3  vss   0.173f
C7  sig7  vss   0.407f
.ends
