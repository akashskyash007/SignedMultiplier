* Spice description of an2_x2
* Spice driver version 134999461
* Date  4/01/2008 at 18:48:26
* vsxlib 0.13um values
.subckt an2_x2 a b vdd vss z
M1a vdd   a     2z    vdd p  L=0.12U  W=1.375U AS=0.364375P AD=0.364375P PS=3.28U   PD=3.28U
M1b 2z    b     vdd   vdd p  L=0.12U  W=1.375U AS=0.364375P AD=0.364375P PS=3.28U   PD=3.28U
M1z z     2z    vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2a n1    a     vss   vss n  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M2b 2z    b     n1    vss n  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M2z vss   2z    z     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C3  2z    vss   0.900f
C5  a     vss   0.716f
C6  b     vss   0.765f
C1  z     vss   0.705f
.ends
