.subckt nd2v6x4 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from nd2v6x4.ext -        technology: scmos
m00 z   b vdd vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 vdd a z   vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 z   b vdd vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m03 vdd a z   vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m04 w1  b z   vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m05 vss a w1  vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
m06 w2  b z   vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m07 vss a w2  vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0  vdd b   0.060f
C1  vdd z   0.135f
C2  vdd a   0.314f
C3  b   z   0.274f
C4  b   a   0.275f
C5  b   w1  0.005f
C6  z   a   0.115f
C7  z   w1  0.018f
C8  z   w2  0.022f
C9  w2  vss 0.023f
C10 w1  vss 0.025f
C11 a   vss 0.330f
C12 z   vss 0.223f
C13 b   vss 0.326f
.ends
