* Spice description of bf1v0x05
* Spice driver version 134999461
* Date  1/01/2008 at 16:39:22
* wsclib 0.13um values
.subckt bf1v0x05 a vdd vss z
M01 an    a     vdd   vdd p  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
M02 an    a     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 vdd   an    z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M04 vss   an    z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C1  an    vss   0.537f
C4  a     vss   0.474f
C3  z     vss   0.476f
.ends
