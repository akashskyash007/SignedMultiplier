* Spice description of inv_x4
* Spice driver version 134999461
* Date  5/01/2008 at 15:08:12
* sxlib 0.13um values
.subckt inv_x4 i nq vdd vss
Mtr_00001 vss   i     nq    vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00002 nq    i     vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00003 vdd   i     nq    vdd p  L=0.12U  W=1.53U  AS=0.40545P  AD=0.40545P  PS=3.59U   PD=3.59U
Mtr_00004 nq    i     vdd   vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C4  i     vss   1.428f
C1  nq    vss   0.784f
.ends
