* Spice description of rowend_x0
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:13
* vsclib 0.13um values
.subckt rowend_x0 vdd vss
.ends
