.subckt nr2av0x4 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2av0x4.ext -        technology: scmos
m00 w1  an vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.428993p ps=2.72907u
m01 z   b  w1  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.19635p  ps=1.795u  
m02 w2  b  z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m03 vdd an w2  vdd p w=1.54u  l=0.13u ad=0.428993p pd=2.72907u as=0.19635p  ps=1.795u  
m04 w3  an vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.428993p ps=2.72907u
m05 z   b  w3  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.19635p  ps=1.795u  
m06 w4  b  z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m07 vdd an w4  vdd p w=1.54u  l=0.13u ad=0.428993p pd=2.72907u as=0.19635p  ps=1.795u  
m08 an  a  vdd vdd p w=1.045u l=0.13u ad=0.21945p  pd=1.465u   as=0.291102p ps=1.85187u
m09 vdd a  an  vdd p w=1.045u l=0.13u ad=0.291102p pd=1.85187u as=0.21945p  ps=1.465u  
m10 z   b  vss vss n w=1.045u l=0.13u ad=0.21945p  pd=1.577u   as=0.418794p ps=2.83316u
m11 vss an z   vss n w=1.045u l=0.13u ad=0.418794p pd=2.83316u as=0.21945p  ps=1.577u  
m12 z   an vss vss n w=0.605u l=0.13u ad=0.12705p  pd=0.913u   as=0.24246p  ps=1.64025u
m13 vss b  z   vss n w=0.605u l=0.13u ad=0.24246p  pd=1.64025u as=0.12705p  ps=0.913u  
m14 vss a  an  vss n w=1.045u l=0.13u ad=0.418794p pd=2.83316u as=0.355575p ps=2.84u   
C0  z   w2  0.009f
C1  an  a   0.090f
C2  z   w3  0.009f
C3  vdd an  0.064f
C4  z   w4  0.004f
C5  vdd b   0.028f
C6  vdd w1  0.004f
C7  vdd z   0.122f
C8  an  b   0.659f
C9  an  w1  0.004f
C10 vdd w2  0.004f
C11 an  z   0.217f
C12 vdd w3  0.004f
C13 an  w2  0.008f
C14 b   z   0.174f
C15 vdd w4  0.004f
C16 vdd a   0.012f
C17 w1  z   0.009f
C18 a   vss 0.143f
C19 w4  vss 0.011f
C20 w3  vss 0.007f
C21 w2  vss 0.007f
C22 z   vss 0.485f
C23 w1  vss 0.008f
C24 b   vss 0.278f
C25 an  vss 0.389f
.ends
