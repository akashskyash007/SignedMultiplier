* Spice description of no2_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:18:30
* ssxlib 0.13um values
.subckt no2_x1 i0 i1 nq vdd vss
Mtr_00001 nq    i0    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00002 vss   i1    nq    vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00003 sig5  i1    nq    vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00004 vdd   i0    sig5  vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
C4  i0    vss   0.981f
C3  i1    vss   0.857f
C1  nq    vss   0.790f
.ends
