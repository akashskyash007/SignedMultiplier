* Spice description of rowend_x0
* Spice driver version 134999461
* Date  4/01/2008 at 19:49:29
* vxlib 0.13um values
.subckt rowend_x0 vdd vss
.ends
