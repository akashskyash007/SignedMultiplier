* Spice description of nd2a_x2
* Spice driver version 134999461
* Date  4/01/2008 at 19:02:55
* vsxlib 0.13um values
.subckt nd2a_x2 a b vdd vss z
M1a 4     a     vdd   vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
M1  z     b     vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2a vss   a     4     vss n  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M2  vdd   4     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3  z     b     sig2  vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
M4  sig2  4     vss   vss n  L=0.12U  W=1.815U AS=0.480975P AD=0.480975P PS=4.16U   PD=4.16U
C5  4     vss   0.815f
C6  a     vss   0.767f
C4  b     vss   0.677f
C1  z     vss   0.797f
.ends
