.subckt buf_x2 i q vdd vss
*05-JAN-08 SPICE3       file   created      from buf_x2.ext -        technology: scmos
m00 vdd i  w1  vdd p w=0.66u  l=0.13u ad=0.230418p pd=1.25882u as=0.2838p   ps=2.18u   
m01 q   w1 vdd vdd p w=2.145u l=0.13u ad=0.92235p  pd=5.15u    as=0.748857p ps=4.09118u
m02 vss i  w1  vss n w=0.33u  l=0.13u ad=0.113586p pd=0.756u   as=0.16005p  ps=1.63u   
m03 q   w1 vss vss n w=1.045u l=0.13u ad=0.44935p  pd=2.95u    as=0.359689p ps=2.394u  
C0 i   q   0.171f
C1 vdd w1  0.010f
C2 vdd i   0.069f
C3 vdd q   0.026f
C4 w1  i   0.184f
C5 q   vss 0.129f
C6 i   vss 0.183f
C7 w1  vss 0.275f
.ends
