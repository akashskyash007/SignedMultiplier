.subckt nd2v4x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v4x1.ext -        technology: scmos
m00 z   b vdd vdd p w=0.99u l=0.13u ad=0.2079p  pd=1.41u  as=0.44385p ps=2.95u 
m01 vdd a z   vdd p w=0.99u l=0.13u ad=0.44385p pd=2.95u  as=0.2079p  ps=1.41u 
m02 w1  b z   vss n w=0.44u l=0.13u ad=0.0561p  pd=0.695u as=0.1529p  ps=1.63u 
m03 vss a w1  vss n w=0.44u l=0.13u ad=0.2981p  pd=2.29u  as=0.0561p  ps=0.695u
C0 b   a   0.108f
C1 b   z   0.085f
C2 a   z   0.009f
C3 a   w1  0.005f
C4 vdd b   0.002f
C5 vdd z   0.086f
C6 w1  vss 0.003f
C7 z   vss 0.162f
C8 a   vss 0.158f
C9 b   vss 0.083f
.ends
