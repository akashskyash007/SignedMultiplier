.subckt aoi22_x2 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from aoi22_x2.ext -        technology: scmos
m00 z   b2 n3  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.561963p ps=3.15625u
m01 n3  b1 z   vdd p w=2.035u l=0.13u ad=0.561963p pd=3.15625u as=0.539275p ps=2.565u  
m02 z   b1 n3  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.561963p ps=3.15625u
m03 n3  b2 z   vdd p w=2.035u l=0.13u ad=0.561963p pd=3.15625u as=0.539275p ps=2.565u  
m04 vdd a2 n3  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.561963p ps=3.15625u
m05 n3  a1 vdd vdd p w=2.035u l=0.13u ad=0.561963p pd=3.15625u as=0.539275p ps=2.565u  
m06 vdd a1 n3  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.561963p ps=3.15625u
m07 n3  a2 vdd vdd p w=2.035u l=0.13u ad=0.561963p pd=3.15625u as=0.539275p ps=2.565u  
m08 w1  b1 vss vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.880275p ps=4.6u    
m09 z   b2 w1  vss n w=1.815u l=0.13u ad=0.480975p pd=2.345u   as=0.281325p ps=2.125u  
m10 w2  a2 z   vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.480975p ps=2.345u  
m11 vss a1 w2  vss n w=1.815u l=0.13u ad=0.880275p pd=4.6u     as=0.281325p ps=2.125u  
C0  z  w1  0.012f
C1  b2 a2  0.161f
C2  b2 n3  0.046f
C3  b2 z   0.220f
C4  b1 n3  0.013f
C5  a2 a1  0.282f
C6  a2 n3  0.155f
C7  b1 z   0.044f
C8  b2 vdd 0.021f
C9  a1 n3  0.013f
C10 b1 vdd 0.021f
C11 b1 w1  0.009f
C12 a2 vdd 0.057f
C13 n3 z   0.204f
C14 a1 vdd 0.021f
C15 n3 vdd 0.308f
C16 z  vdd 0.030f
C17 b2 b1  0.282f
C18 w2 vss 0.020f
C19 w1 vss 0.016f
C21 z  vss 0.413f
C22 n3 vss 0.171f
C23 a1 vss 0.158f
C24 a2 vss 0.208f
C25 b1 vss 0.139f
C26 b2 vss 0.212f
.ends
