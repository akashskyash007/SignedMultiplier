.subckt mxn2v2x1 a0 a1 s vdd vss z
*01-JAN-08 SPICE3       file   created      from mxn2v2x1.ext -        technology: scmos
m00 vdd a0  a0n vdd p w=0.715u l=0.13u ad=0.245513p pd=1.64613u as=0.225775p ps=2.18u   
m01 a0i a0n vdd vdd p w=1.21u  l=0.13u ad=0.2541p   pd=1.63u    as=0.415484p ps=2.78575u
m02 z   s   a0i vdd p w=1.21u  l=0.13u ad=0.2541p   pd=1.63u    as=0.2541p   ps=1.63u   
m03 a1i sn  z   vdd p w=1.21u  l=0.13u ad=0.3872p   pd=1.85u    as=0.2541p   ps=1.63u   
m04 vdd a1n a1i vdd p w=1.21u  l=0.13u ad=0.415484p pd=2.78575u as=0.3872p   ps=1.85u   
m05 vdd a1  a1n vdd p w=0.715u l=0.13u ad=0.245513p pd=1.64613u as=0.225775p ps=2.18u   
m06 sn  s   vdd vdd p w=0.55u  l=0.13u ad=0.18205p  pd=1.85u    as=0.188856p ps=1.26625u
m07 vss a0  a0n vss n w=0.55u  l=0.13u ad=0.192051p pd=1.46122u as=0.18205p  ps=1.85u   
m08 a0i a0n vss vss n w=0.605u l=0.13u ad=0.12705p  pd=1.025u   as=0.211256p ps=1.60735u
m09 z   sn  a0i vss n w=0.605u l=0.13u ad=0.142175p pd=1.3u     as=0.12705p  ps=1.025u  
m10 a1i s   z   vss n w=0.605u l=0.13u ad=0.136125p pd=1.19u    as=0.142175p ps=1.3u    
m11 vss a1n a1i vss n w=0.605u l=0.13u ad=0.211256p pd=1.60735u as=0.136125p ps=1.19u   
m12 vss a1  a1n vss n w=0.55u  l=0.13u ad=0.192051p pd=1.46122u as=0.18205p  ps=1.85u   
m13 sn  s   vss vss n w=0.385u l=0.13u ad=0.144375p pd=1.52u    as=0.134436p ps=1.02286u
C0  s   sn  0.125f
C1  z   a1i 0.051f
C2  a0n sn  0.027f
C3  s   a1n 0.029f
C4  vdd z   0.043f
C5  a0n a0  0.164f
C6  sn  a1n 0.080f
C7  vdd a1  0.014f
C8  a0n a0i 0.109f
C9  s   z   0.007f
C10 a0n z   0.027f
C11 sn  a0i 0.028f
C12 sn  z   0.120f
C13 s   a1  0.094f
C14 vdd s   0.062f
C15 sn  a1i 0.107f
C16 vdd a0n 0.050f
C17 a1n a1i 0.015f
C18 sn  a1  0.072f
C19 vdd sn  0.068f
C20 a0i z   0.139f
C21 a1n a1  0.055f
C22 vdd a1n 0.002f
C23 s   a0n 0.040f
C24 a1  vss 0.087f
C25 a1i vss 0.078f
C26 z   vss 0.078f
C27 a0i vss 0.050f
C28 a0  vss 0.124f
C29 a1n vss 0.146f
C30 sn  vss 0.210f
C31 a0n vss 0.170f
C32 s   vss 0.413f
.ends
