.subckt an2v0x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from an2v0x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.41965p   pd=2.86788u as=0.48675p   ps=3.83u   
m01 zn  a  vdd vdd p w=1.045u l=0.13u ad=0.21945p   pd=1.465u   as=0.284763p  ps=1.94606u
m02 vdd b  zn  vdd p w=1.045u l=0.13u ad=0.284763p  pd=1.94606u as=0.21945p   ps=1.465u  
m03 vss zn z   vss n w=0.77u  l=0.13u ad=0.329532p  pd=1.91852u as=0.28875p   ps=2.29u   
m04 w1  a  vss vss n w=0.715u l=0.13u ad=0.0911625p pd=0.97u    as=0.305994p  ps=1.78148u
m05 zn  b  w1  vss n w=0.715u l=0.13u ad=0.225775p  pd=2.18u    as=0.0911625p ps=0.97u   
C0  zn a   0.160f
C1  zn b   0.036f
C2  zn z   0.137f
C3  a  b   0.151f
C4  a  z   0.006f
C5  zn vdd 0.092f
C6  a  vdd 0.007f
C7  zn w1  0.008f
C8  b  vdd 0.032f
C9  a  w1  0.007f
C10 z  vdd 0.034f
C11 w1 vss 0.003f
C13 z  vss 0.228f
C14 b  vss 0.095f
C15 a  vss 0.099f
C16 zn vss 0.211f
.ends
