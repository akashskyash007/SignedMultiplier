.subckt vfeed3 vdd vss
*04-JAN-08 SPICE3       file   created      from vfeed3.ext -        technology: scmos
.ends
