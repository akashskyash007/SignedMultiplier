* Spice description of bf1v5x05
* Spice driver version 134999461
* Date  1/01/2008 at 16:40:57
* vsclib 0.13um values
.subckt bf1v5x05 a vdd vss z
M01 an    a     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M02 an    a     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M03 vdd   an    z     vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M04 vss   an    z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C2  an    vss   0.407f
C4  a     vss   0.457f
C3  z     vss   0.485f
.ends
