.subckt ao22_x4 i0 i1 i2 q vdd vss
*05-JAN-08 SPICE3       file   created      from ao22_x4.ext -        technology: scmos
m00 w1  i0 vdd vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.6718u  as=0.556059p ps=2.55932u
m01 w2  i1 w1  vdd p w=1.045u l=0.13u ad=0.276925p pd=1.58821u as=0.276925p ps=1.58821u
m02 vdd i2 w2  vdd p w=1.1u   l=0.13u ad=0.556059p pd=2.55932u as=0.2915p   ps=1.6718u 
m03 q   w2 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=1.08432p  ps=4.99068u
m04 vdd w2 q   vdd p w=2.145u l=0.13u ad=1.08432p  pd=4.99068u as=0.568425p ps=2.675u  
m05 w2  i0 w3  vss n w=0.55u  l=0.13u ad=0.21835p  pd=1.52u    as=0.177043p ps=1.42069u
m06 w3  i1 w2  vss n w=0.55u  l=0.13u ad=0.177043p pd=1.42069u as=0.21835p  ps=1.52u   
m07 vss i2 w3  vss n w=0.495u l=0.13u ad=0.244709p pd=1.29447u as=0.159339p ps=1.27862u
m08 q   w2 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.516608p ps=2.73277u
m09 vss w2 q   vss n w=1.045u l=0.13u ad=0.516608p pd=2.73277u as=0.276925p ps=1.575u  
C0  w2  q   0.007f
C1  i1  i2  0.051f
C2  w2  w3  0.062f
C3  i1  w1  0.034f
C4  i0  w3  0.007f
C5  i1  w3  0.007f
C6  vdd w2  0.033f
C7  i2  w3  0.012f
C8  vdd i0  0.037f
C9  vdd i1  0.015f
C10 vdd i2  0.062f
C11 w2  i1  0.145f
C12 vdd q   0.080f
C13 w2  i2  0.192f
C14 i0  i1  0.207f
C15 w3  vss 0.125f
C16 q   vss 0.136f
C17 w1  vss 0.008f
C18 i2  vss 0.184f
C19 i1  vss 0.144f
C20 i0  vss 0.149f
C21 w2  vss 0.322f
.ends
