* Spice description of inv_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:08:08
* ssxlib 0.13um values
.subckt inv_x2 i nq vdd vss
Mtr_00001 vss   i     nq    vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 nq    i     vdd   vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
C3  i     vss   0.914f
C1  nq    vss   0.714f
.ends
