.subckt oa2a22_x4 i0 i1 i2 i3 q vdd vss
*05-JAN-08 SPICE3       file   created      from oa2a22_x4.ext -        technology: scmos
m00 w1  i0 w2  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.38225p  ps=2.345u  
m01 w2  i1 w1  vdd p w=1.1u   l=0.13u ad=0.38225p  pd=2.345u   as=0.2915p   ps=1.63u   
m02 vdd i2 w2  vdd p w=1.1u   l=0.13u ad=0.436085p pd=2.44746u as=0.38225p  ps=2.345u  
m03 w2  i3 vdd vdd p w=1.1u   l=0.13u ad=0.38225p  pd=2.345u   as=0.436085p ps=2.44746u
m04 q   w1 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.850365p ps=4.77254u
m05 vdd w1 q   vdd p w=2.145u l=0.13u ad=0.850365p pd=4.77254u as=0.568425p ps=2.675u  
m06 w3  i0 vss vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.286569p ps=1.99655u
m07 w1  i1 w3  vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.14575p  ps=1.08u   
m08 w4  i2 w1  vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.14575p  ps=1.08u   
m09 vss i3 w4  vss n w=0.55u  l=0.13u ad=0.286569p pd=1.99655u as=0.14575p  ps=1.08u   
m10 q   w1 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.544481p ps=3.79345u
m11 vss w1 q   vss n w=1.045u l=0.13u ad=0.544481p pd=3.79345u as=0.276925p ps=1.575u  
C0  w1  i2  0.138f
C1  vdd w2  0.165f
C2  i0  i1  0.208f
C3  w1  i3  0.019f
C4  vdd q   0.092f
C5  w1  w2  0.163f
C6  i1  i2  0.078f
C7  w1  q   0.098f
C8  i0  w2  0.007f
C9  i1  w2  0.007f
C10 i2  i3  0.208f
C11 i2  w2  0.007f
C12 vdd w1  0.088f
C13 i1  w3  0.017f
C14 i3  w2  0.007f
C15 vdd i0  0.003f
C16 vdd i1  0.003f
C17 i2  w4  0.017f
C18 vdd i2  0.003f
C19 w1  i1  0.138f
C20 vdd i3  0.003f
C21 w4  vss 0.005f
C22 w3  vss 0.005f
C23 q   vss 0.147f
C24 w2  vss 0.084f
C25 i3  vss 0.178f
C26 i2  vss 0.178f
C27 i1  vss 0.178f
C28 i0  vss 0.179f
C29 w1  vss 0.354f
.ends
