.subckt aoi211v0x05 a1 a2 b c vdd vss z
*01-JAN-08 SPICE3       file   created      from aoi211v0x05.ext -        technology: scmos
m00 w1  c  z   vdd p w=1.54u  l=0.13u ad=0.19635p   pd=1.795u    as=0.48675p   ps=3.83u    
m01 n1  b  w1  vdd p w=1.54u  l=0.13u ad=0.363733p  pd=2.58333u  as=0.19635p   ps=1.795u   
m02 vdd a1 n1  vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u     as=0.363733p  ps=2.58333u 
m03 n1  a2 vdd vdd p w=1.54u  l=0.13u ad=0.363733p  pd=2.58333u  as=0.3234p    ps=1.96u    
m04 z   c  vss vss n w=0.33u  l=0.13u ad=0.08745p   pd=0.925714u as=0.219686p  ps=1.80571u 
m05 vss b  z   vss n w=0.33u  l=0.13u ad=0.219686p  pd=1.80571u  as=0.08745p   ps=0.925714u
m06 w2  a1 vss vss n w=0.495u l=0.13u ad=0.0631125p pd=0.75u     as=0.329529p  ps=2.70857u 
m07 z   a2 w2  vss n w=0.495u l=0.13u ad=0.131175p  pd=1.38857u  as=0.0631125p ps=0.75u    
C0  z  w2  0.009f
C1  w1 vdd 0.004f
C2  n1 vdd 0.098f
C3  b  a1  0.103f
C4  b  a2  0.023f
C5  c  z   0.146f
C6  b  z   0.100f
C7  a1 a2  0.134f
C8  a1 z   0.057f
C9  a2 z   0.007f
C10 b  n1  0.070f
C11 c  vdd 0.007f
C12 a1 n1  0.006f
C13 b  vdd 0.012f
C14 z  w1  0.005f
C15 a2 n1  0.080f
C16 a1 vdd 0.007f
C17 a2 vdd 0.019f
C18 z  vdd 0.017f
C19 c  b   0.110f
C20 w2 vss 0.004f
C22 n1 vss 0.020f
C23 w1 vss 0.009f
C24 z  vss 0.235f
C25 a2 vss 0.131f
C26 a1 vss 0.097f
C27 b  vss 0.094f
C28 c  vss 0.211f
.ends
