* Spice description of or2v0x2
* Spice driver version 134999461
* Date  1/01/2008 at 17:00:17
* wsclib 0.13um values
.subckt or2v0x2 a b vdd vss z
M01 03    a     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 sig1  a     vss   vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M03 sig1  b     03    vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 vss   b     sig1  vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
M05 vdd   sig1  z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M06 vss   sig1  z     vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C4  a     vss   0.441f
C5  b     vss   0.658f
C1  sig1  vss   0.638f
C2  z     vss   0.703f
.ends
