.subckt dfnt1v0x2 cp d vdd vss z
*01-JAN-08 SPICE3       file   created      from dfnt1v0x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.409794p  pd=3.3124u   as=0.4928p    ps=3.83u   
m01 zn  n4 vdd vdd p w=0.77u  l=0.13u ad=0.24035p   pd=2.29u     as=0.204897p  ps=1.6562u 
m02 w1  zn vdd vdd p w=0.33u  l=0.13u ad=0.042075p  pd=0.585u    as=0.087813p  ps=0.7098u 
m03 n4  ci w1  vdd p w=0.33u  l=0.13u ad=0.07535p   pd=0.72u     as=0.042075p  ps=0.585u  
m04 n2  cn n4  vdd p w=0.66u  l=0.13u ad=0.1386p    pd=1.08u     as=0.1507p    ps=1.44u   
m05 vdd n1 n2  vdd p w=0.66u  l=0.13u ad=0.175626p  pd=1.4196u   as=0.1386p    ps=1.08u   
m06 w2  n2 vdd vdd p w=0.33u  l=0.13u ad=0.042075p  pd=0.585u    as=0.087813p  ps=0.7098u 
m07 n1  cn w2  vdd p w=0.33u  l=0.13u ad=0.0759868p pd=0.716842u as=0.042075p  ps=0.585u  
m08 vss zn z   vss n w=0.77u  l=0.13u ad=0.223765p  pd=2.21828u  as=0.24035p   ps=2.29u   
m09 vss n4 zn  vss n w=0.385u l=0.13u ad=0.111882p  pd=1.10914u  as=0.138325p  ps=1.52u   
m10 w3  ci n1  vdd p w=0.715u l=0.13u ad=0.0911625p pd=0.97u     as=0.164638p  ps=1.55316u
m11 vdd d  w3  vdd p w=0.715u l=0.13u ad=0.190262p  pd=1.5379u   as=0.0911625p ps=0.97u   
m12 ci  cn vdd vdd p w=0.605u l=0.13u ad=0.196625p  pd=1.96u     as=0.160991p  ps=1.3013u 
m13 cn  cp vdd vdd p w=0.55u  l=0.13u ad=0.18205p   pd=1.85u     as=0.146355p  ps=1.183u  
m14 vss cn ci  vss n w=0.33u  l=0.13u ad=0.0958992p pd=0.95069u  as=0.12375p   ps=1.41u   
m15 w4  zn vss vss n w=0.33u  l=0.13u ad=0.042075p  pd=0.585u    as=0.0958992p ps=0.95069u
m16 n4  cn w4  vss n w=0.33u  l=0.13u ad=0.0693p    pd=0.75u     as=0.042075p  ps=0.585u  
m17 n2  ci n4  vss n w=0.33u  l=0.13u ad=0.0693p    pd=0.75u     as=0.0693p    ps=0.75u   
m18 vss n1 n2  vss n w=0.33u  l=0.13u ad=0.0958992p pd=0.95069u  as=0.0693p    ps=0.75u   
m19 w5  n2 vss vss n w=0.33u  l=0.13u ad=0.042075p  pd=0.585u    as=0.0958992p ps=0.95069u
m20 n1  ci w5  vss n w=0.33u  l=0.13u ad=0.0693p    pd=0.75u     as=0.042075p  ps=0.585u  
m21 w6  cn n1  vss n w=0.33u  l=0.13u ad=0.042075p  pd=0.585u    as=0.0693p    ps=0.75u   
m22 vss d  w6  vss n w=0.33u  l=0.13u ad=0.0958992p pd=0.95069u  as=0.042075p  ps=0.585u  
m23 cn  cp vss vss n w=0.385u l=0.13u ad=0.144375p  pd=1.52u     as=0.111882p  ps=1.10914u
C0  cp  cn  0.128f
C1  vdd z   0.030f
C2  ci  cn  0.246f
C3  vdd cn  0.074f
C4  ci  n4  0.090f
C5  ci  n1  0.179f
C6  n4  w4  0.010f
C7  n4  vdd 0.041f
C8  zn  z   0.050f
C9  vdd n1  0.043f
C10 d   cp  0.006f
C11 ci  n2  0.120f
C12 w5  n1  0.008f
C13 ci  d   0.190f
C14 vdd n2  0.012f
C15 zn  cn  0.055f
C16 d   vdd 0.003f
C17 n4  zn  0.116f
C18 ci  w3  0.005f
C19 ci  cp  0.027f
C20 cp  vdd 0.023f
C21 n4  cn  0.011f
C22 cn  n1  0.076f
C23 ci  vdd 0.039f
C24 cn  n2  0.073f
C25 d   cn  0.105f
C26 n4  w1  0.008f
C27 n4  n2  0.019f
C28 n1  n2  0.167f
C29 ci  zn  0.050f
C30 w2  n1  0.003f
C31 vdd zn  0.007f
C32 w6  vss 0.004f
C33 w5  vss 0.002f
C34 w4  vss 0.002f
C35 cp  vss 0.114f
C36 w3  vss 0.004f
C37 w2  vss 0.001f
C38 n4  vss 0.213f
C39 d   vss 0.119f
C40 ci  vss 0.377f
C41 n2  vss 0.184f
C42 n1  vss 0.247f
C43 cn  vss 0.439f
C44 z   vss 0.142f
C45 zn  vss 0.251f
.ends
