.subckt nr2av0x1 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from nr2av0x1.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.43u l=0.13u ad=0.431383p pd=2.51u  as=0.53625p  ps=3.61u 
m01 w2  a   vdd vdd p w=1.43u l=0.13u ad=0.53625p  pd=3.61u  as=0.431383p ps=2.51u 
m02 w3  w2  vdd vdd p w=1.43u l=0.13u ad=0.37895p  pd=1.96u  as=0.431383p ps=2.51u 
m03 z   b   w3  vdd p w=1.43u l=0.13u ad=0.53625p  pd=3.61u  as=0.37895p  ps=1.96u 
m04 vss vss w4  vss n w=0.99u l=0.13u ad=0.3168p   pd=2.125u as=0.37125p  ps=2.73u 
m05 w2  a   vss vss n w=0.99u l=0.13u ad=0.37125p  pd=2.73u  as=0.3168p   ps=2.125u
m06 z   w2  vss vss n w=0.99u l=0.13u ad=0.26235p  pd=1.52u  as=0.3168p   ps=2.125u
m07 vss b   z   vss n w=0.99u l=0.13u ad=0.3168p   pd=2.125u as=0.26235p  ps=1.52u 
C0  w2  b   0.129f
C1  w2  z   0.089f
C2  b   z   0.144f
C3  vdd a   0.100f
C4  w3  z   0.020f
C5  vdd w2  0.059f
C6  vdd b   0.009f
C7  a   w2  0.093f
C8  w4  vss 0.011f
C9  z   vss 0.106f
C10 w3  vss 0.014f
C11 w1  vss 0.014f
C12 b   vss 0.215f
C13 w2  vss 0.334f
C14 a   vss 0.291f
.ends
