.subckt fulladder_x4 a1 a2 a3 a4 b1 b2 b3 b4 cin1 cin2 cin3 cout sout vdd vss
*05-JAN-08 SPICE3       file   created      from fulladder_x4.ext -        technology: scmos
m00 vdd  a1   w1   vdd p w=0.98u l=0.13u ad=0.335205p pd=1.83562u  as=0.346012p ps=2.13982u 
m01 w1   b1   vdd  vdd p w=0.98u l=0.13u ad=0.346012p pd=2.13982u  as=0.335205p ps=1.83562u 
m02 w2   cin1 w1   vdd p w=0.98u l=0.13u ad=0.278565p pd=1.5925u   as=0.346012p ps=2.13982u 
m03 w3   a2   w2   vdd p w=1.42u l=0.13u ad=0.2982p   pd=1.84u     as=0.403635p ps=2.3075u  
m04 w1   b2   w3   vdd p w=1.42u l=0.13u ad=0.501364p pd=3.10055u  as=0.2982p   ps=1.84u    
m05 w4   a1   vss  vss n w=0.54u l=0.13u ad=0.11315p  pd=0.971092u as=0.217718p ps=1.49655u 
m06 w2   b1   w4   vss n w=0.65u l=0.13u ad=0.193435p pd=1.42037u  as=0.1362p   ps=1.16891u 
m07 cout w2   vdd  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u     as=0.749081p ps=4.10204u 
m08 vdd  w2   cout vdd p w=2.19u l=0.13u ad=0.749081p pd=4.10204u  as=0.58035p  ps=2.72u    
m09 sout w5   vdd  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u     as=0.749081p ps=4.10204u 
m10 vdd  w5   sout vdd p w=2.19u l=0.13u ad=0.749081p pd=4.10204u  as=0.58035p  ps=2.72u    
m11 w6   a3   vdd  vdd p w=0.76u l=0.13u ad=0.244353p pd=1.58995u  as=0.259955p ps=1.42354u 
m12 vdd  b3   w6   vdd p w=0.76u l=0.13u ad=0.259955p pd=1.42354u  as=0.244353p ps=1.58995u 
m13 w6   cin2 vdd  vdd p w=0.76u l=0.13u ad=0.244353p pd=1.58995u  as=0.259955p ps=1.42354u 
m14 w5   w2   w6   vdd p w=0.98u l=0.13u ad=0.27271p  pd=1.70092u  as=0.315087p ps=2.0502u  
m15 w7   cin3 w5   vdd p w=0.76u l=0.13u ad=0.1596p   pd=1.18u     as=0.21149p  ps=1.31908u 
m16 w8   a4   w7   vdd p w=0.76u l=0.13u ad=0.1596p   pd=1.18u     as=0.1596p   ps=1.18u    
m17 w6   b4   w8   vdd p w=0.76u l=0.13u ad=0.244353p pd=1.58995u  as=0.1596p   ps=1.18u    
m18 w9   cin1 w2   vss n w=0.43u l=0.13u ad=0.136883p pd=1.21u     as=0.127965p ps=0.93963u 
m19 vss  a2   w9   vss n w=0.43u l=0.13u ad=0.173368p pd=1.1917u   as=0.136883p ps=1.21u    
m20 w9   b2   vss  vss n w=0.43u l=0.13u ad=0.136883p pd=1.21u     as=0.173368p ps=1.1917u  
m21 cout w2   vss  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u     as=0.439468p ps=3.02082u 
m22 vss  w2   cout vss n w=1.09u l=0.13u ad=0.439468p pd=3.02082u  as=0.28885p  ps=1.62u    
m23 sout w5   vss  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u     as=0.439468p ps=3.02082u 
m24 vss  w5   sout vss n w=1.09u l=0.13u ad=0.439468p pd=3.02082u  as=0.28885p  ps=1.62u    
m25 w10  a3   vss  vss n w=0.43u l=0.13u ad=0.0903p   pd=0.85u     as=0.173368p ps=1.1917u  
m26 w11  b3   w10  vss n w=0.43u l=0.13u ad=0.0903p   pd=0.85u     as=0.0903p   ps=0.85u    
m27 w5   cin2 w11  vss n w=0.43u l=0.13u ad=0.111024p pd=0.94866u  as=0.0903p   ps=0.85u    
m28 w12  w2   w5   vss n w=0.54u l=0.13u ad=0.141152p pd=1.19803u  as=0.139426p ps=1.19134u 
m29 vss  cin3 w12  vss n w=0.43u l=0.13u ad=0.173368p pd=1.1917u   as=0.112399p ps=0.953989u
m30 w12  a4   vss  vss n w=0.43u l=0.13u ad=0.112399p pd=0.953989u as=0.173368p ps=1.1917u  
m31 vss  b4   w12  vss n w=0.43u l=0.13u ad=0.173368p pd=1.1917u   as=0.112399p ps=0.953989u
C0  b2   w9   0.014f
C1  b3   cin2 0.189f
C2  w5   cin3 0.073f
C3  w2   w1   0.119f
C4  b1   cin1 0.073f
C5  b3   w6   0.005f
C6  w2   w3   0.011f
C7  vdd  w6   0.171f
C8  cin2 w6   0.005f
C9  a1   w1   0.023f
C10 cin1 a2   0.162f
C11 cin3 w12  0.014f
C12 w2   cout 0.100f
C13 b1   w1   0.014f
C14 vdd  w1   0.156f
C15 a4   w12  0.015f
C16 w6   cin3 0.006f
C17 w2   w9   0.009f
C18 w2   sout 0.034f
C19 cin1 w1   0.005f
C20 a2   b2   0.182f
C21 w2   w5   0.184f
C22 w6   a4   0.014f
C23 w5   sout 0.050f
C24 w2   a3   0.014f
C25 b1   w4   0.002f
C26 a2   w1   0.005f
C27 w6   b4   0.023f
C28 cin3 a4   0.179f
C29 w5   w10  0.011f
C30 w2   b3   0.014f
C31 a2   w3   0.007f
C32 b2   w1   0.012f
C33 w5   a3   0.085f
C34 w2   b1   0.095f
C35 vdd  cout 0.019f
C36 vdd  w2   0.221f
C37 w5   w11  0.011f
C38 w5   b3   0.021f
C39 w2   cin2 0.145f
C40 w2   cin1 0.096f
C41 vdd  sout 0.019f
C42 vdd  w5   0.020f
C43 a4   b4   0.206f
C44 w5   w12  0.016f
C45 cin1 w9   0.010f
C46 a3   b3   0.157f
C47 w5   cin2 0.021f
C48 w2   w6   0.077f
C49 w1   w3   0.011f
C50 w2   a2   0.014f
C51 a1   b1   0.200f
C52 a2   w9   0.014f
C53 w5   w6   0.021f
C54 w2   cin3 0.061f
C55 w2   b2   0.014f
C56 vdd  b1   0.015f
C57 a4   w8   0.009f
C58 w12  vss  0.110f
C59 w11  vss  0.006f
C60 w10  vss  0.005f
C61 w9   vss  0.114f
C62 w8   vss  0.006f
C63 w7   vss  0.006f
C64 b4   vss  0.133f
C65 a4   vss  0.143f
C66 cin3 vss  0.138f
C67 w6   vss  0.076f
C68 cin2 vss  0.142f
C69 b3   vss  0.135f
C70 a3   vss  0.132f
C71 sout vss  0.129f
C72 cout vss  0.137f
C73 w4   vss  0.007f
C74 w3   vss  0.015f
C75 w1   vss  0.072f
C76 b2   vss  0.112f
C77 a2   vss  0.127f
C78 cin1 vss  0.146f
C79 b1   vss  0.142f
C80 a1   vss  0.169f
C81 w5   vss  0.383f
C82 w2   vss  0.481f
.ends
