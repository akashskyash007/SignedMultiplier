.subckt noa2a2a2a24_x4 i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa2a2a2a24_x4.ext -        technology: scmos
m00 w1  i7 w2  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.726275p ps=3.83u   
m01 w2  i6 w1  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.55385p  ps=2.62u   
m02 w2  i5 w3  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.726275p ps=3.83u   
m03 w3  i4 w2  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.726275p ps=3.83u   
m04 w4  i3 w3  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.61312u as=0.726275p ps=3.83u   
m05 w3  i2 w4  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.55385p  ps=2.61312u
m06 w4  i1 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.68188u as=0.685059p ps=3.51222u
m07 vdd i0 w4  vdd p w=2.145u l=0.13u ad=0.685059p pd=3.51222u as=0.568425p ps=2.68188u
m08 nq  w5 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.685059p ps=3.51222u
m09 vdd w5 nq  vdd p w=2.145u l=0.13u ad=0.685059p pd=3.51222u as=0.568425p ps=2.675u  
m10 w5  w1 vdd vdd p w=1.1u   l=0.13u ad=0.473p    pd=3.06u    as=0.351313p ps=1.80114u
m11 w6  i7 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.368044p ps=2.34024u
m12 w1  i6 w6  vss n w=1.045u l=0.13u ad=0.361988p pd=2.2648u  as=0.276925p ps=1.575u  
m13 w7  i5 vss vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.368044p ps=2.34024u
m14 w1  i4 w7  vss n w=1.045u l=0.13u ad=0.361988p pd=2.2648u  as=0.161975p ps=1.355u  
m15 w8  i3 w1  vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.361988p ps=2.2648u 
m16 vss i2 w8  vss n w=1.045u l=0.13u ad=0.368044p pd=2.34024u as=0.161975p ps=1.355u  
m17 w9  i1 w1  vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.342936p ps=2.1456u 
m18 vss i0 w9  vss n w=0.99u  l=0.13u ad=0.348673p pd=2.21707u as=0.15345p  ps=1.3u    
m19 nq  w5 vss vss n w=1.045u l=0.13u ad=0.349525p pd=2.015u   as=0.368044p ps=2.34024u
m20 vss w5 nq  vss n w=1.045u l=0.13u ad=0.368044p pd=2.34024u as=0.349525p ps=2.015u  
m21 w5  w1 vss vss n w=0.55u  l=0.13u ad=0.2365p   pd=1.96u    as=0.193707p ps=1.23171u
C0  i3  vdd 0.010f
C1  vdd i7  0.010f
C2  w1  w8  0.010f
C3  i5  w1  0.019f
C4  i0  w1  0.019f
C5  i2  w4  0.034f
C6  i4  i3  0.200f
C7  i2  vdd 0.010f
C8  w1  w9  0.010f
C9  i5  w3  0.007f
C10 i1  w4  0.025f
C11 w5  w1  0.159f
C12 i1  vdd 0.016f
C13 i0  w4  0.008f
C14 w2  w1  0.059f
C15 i6  w2  0.037f
C16 i5  vdd 0.010f
C17 i3  i2  0.232f
C18 i0  vdd 0.053f
C19 i5  i4  0.232f
C20 i0  nq  0.119f
C21 w2  w3  0.097f
C22 i6  w1  0.112f
C23 w5  vdd 0.032f
C24 w5  nq  0.020f
C25 w2  vdd 0.122f
C26 i4  w2  0.005f
C27 w1  vdd 0.017f
C28 i6  vdd 0.010f
C29 w1  nq  0.040f
C30 w3  w4  0.088f
C31 i4  w1  0.019f
C32 i1  i0  0.124f
C33 w2  i7  0.016f
C34 w3  vdd 0.192f
C35 i3  w1  0.019f
C36 i4  w3  0.012f
C37 w1  i7  0.117f
C38 w4  vdd 0.097f
C39 i6  i7  0.096f
C40 w1  w6  0.015f
C41 i2  w1  0.019f
C42 i3  w3  0.016f
C43 i0  w5  0.100f
C44 nq  vdd 0.072f
C45 i4  vdd 0.010f
C46 w1  w7  0.010f
C47 i5  w2  0.028f
C48 i1  w1  0.019f
C49 i2  w3  0.007f
C50 w9  vss 0.014f
C51 w8  vss 0.014f
C52 w7  vss 0.014f
C53 w6  vss 0.025f
C54 nq  vss 0.096f
C55 w4  vss 0.066f
C56 w3  vss 0.107f
C57 w1  vss 0.816f
C58 w2  vss 0.125f
C59 w5  vss 0.291f
C60 i0  vss 0.159f
C61 i1  vss 0.134f
C62 i2  vss 0.129f
C63 i3  vss 0.136f
C64 i4  vss 0.124f
C65 i5  vss 0.135f
C66 i6  vss 0.150f
C67 i7  vss 0.169f
.ends
