.subckt inv_x8 i nq vdd vss
*05-JAN-08 SPICE3       file   created      from inv_x8.ext -        technology: scmos
m00 nq  i vdd vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.689p   ps=3.975u
m01 vdd i nq  vdd p w=2.19u l=0.13u ad=0.689p   pd=3.975u as=0.58035p ps=2.72u 
m02 nq  i vdd vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.689p   ps=3.975u
m03 vdd i nq  vdd p w=2.19u l=0.13u ad=0.689p   pd=3.975u as=0.58035p ps=2.72u 
m04 nq  i vss vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.37605p ps=2.325u
m05 vss i nq  vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.28885p ps=1.62u 
m06 nq  i vss vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.37605p ps=2.325u
m07 vss i nq  vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.28885p ps=1.62u 
C0 vdd i   0.103f
C1 vdd nq  0.183f
C2 i   nq  0.220f
C3 nq  vss 0.316f
C4 i   vss 0.486f
.ends
