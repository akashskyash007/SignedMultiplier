.subckt nd3_x2 a b c vdd vss z
*04-JAN-08 SPICE3       file   created      from nd3_x2.ext -        technology: scmos
m00 vdd c z   vdd p w=1.815u l=0.13u ad=0.5808p   pd=3.06u  as=0.523325p ps=3.06u 
m01 z   b vdd vdd p w=1.815u l=0.13u ad=0.523325p pd=3.06u  as=0.5808p   ps=3.06u 
m02 vdd a z   vdd p w=1.815u l=0.13u ad=0.5808p   pd=3.06u  as=0.523325p ps=3.06u 
m03 w1  c z   vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u as=0.535425p ps=4.49u 
m04 w2  b w1  vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u as=0.281325p ps=2.125u
m05 vss a w2  vss n w=1.815u l=0.13u ad=0.78045p  pd=4.49u  as=0.281325p ps=2.125u
C0  c  b   0.193f
C1  c  a   0.066f
C2  c  z   0.094f
C3  b  a   0.201f
C4  b  z   0.059f
C5  c  vdd 0.016f
C6  b  vdd 0.025f
C7  a  z   0.030f
C8  c  w1  0.005f
C9  a  vdd 0.010f
C10 c  w2  0.002f
C11 a  w1  0.012f
C12 z  vdd 0.104f
C13 a  w2  0.012f
C14 w2 vss 0.020f
C15 w1 vss 0.018f
C17 z  vss 0.203f
C18 a  vss 0.119f
C19 b  vss 0.129f
C20 c  vss 0.146f
.ends
