.subckt oa2a22_x2 i0 i1 i2 i3 q vdd vss
*05-JAN-08 SPICE3       file   created      from oa2a22_x2.ext -        technology: scmos
m00 w1  i0 w2  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.38225p  ps=2.345u  
m01 w2  i1 w1  vdd p w=1.1u   l=0.13u ad=0.38225p  pd=2.345u   as=0.2915p   ps=1.63u   
m02 vdd i2 w2  vdd p w=1.1u   l=0.13u ad=0.417861p pd=2.3519u  as=0.38225p  ps=2.345u  
m03 w2  i3 vdd vdd p w=1.1u   l=0.13u ad=0.38225p  pd=2.345u   as=0.417861p ps=2.3519u 
m04 q   w1 vdd vdd p w=2.145u l=0.13u ad=0.92235p  pd=5.15u    as=0.814829p ps=4.5862u 
m05 w3  i0 vss vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.310962p ps=2.21282u
m06 w1  i1 w3  vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.14575p  ps=1.08u   
m07 w4  i2 w1  vss n w=0.55u  l=0.13u ad=0.14575p  pd=1.08u    as=0.14575p  ps=1.08u   
m08 vss i3 w4  vss n w=0.55u  l=0.13u ad=0.310962p pd=2.21282u as=0.14575p  ps=1.08u   
m09 q   w1 vss vss n w=1.045u l=0.13u ad=0.44935p  pd=2.95u    as=0.590827p ps=4.20436u
C0  vdd i3  0.003f
C1  w1  i1  0.138f
C2  vdd w2  0.165f
C3  w1  i2  0.138f
C4  i0  i1  0.208f
C5  w1  i3  0.019f
C6  vdd q   0.038f
C7  w1  w2  0.163f
C8  i1  i2  0.078f
C9  w1  q   0.091f
C10 i0  w2  0.007f
C11 i1  w2  0.007f
C12 i2  i3  0.208f
C13 i2  w2  0.007f
C14 i3  w2  0.007f
C15 vdd w1  0.078f
C16 i1  w3  0.017f
C17 vdd i0  0.003f
C18 vdd i1  0.003f
C19 i2  w4  0.017f
C20 vdd i2  0.003f
C21 w4  vss 0.005f
C22 w3  vss 0.005f
C23 q   vss 0.130f
C24 w2  vss 0.084f
C25 i3  vss 0.178f
C26 i2  vss 0.178f
C27 i1  vss 0.178f
C28 i0  vss 0.179f
C29 w1  vss 0.264f
.ends
