.subckt no3_x4 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from no3_x4.ext -        technology: scmos
m00 w1  i2 w2  vdd p w=2.19u l=0.13u ad=0.33945p  pd=2.5u     as=0.93075p  ps=5.23u   
m01 w3  i1 w1  vdd p w=2.19u l=0.13u ad=0.33945p  pd=2.5u     as=0.33945p  ps=2.5u    
m02 vdd i0 w3  vdd p w=2.19u l=0.13u ad=0.768416p pd=3.2364u  as=0.33945p  ps=2.5u    
m03 nq  w4 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.768416p ps=3.2364u 
m04 vdd w4 nq  vdd p w=2.19u l=0.13u ad=0.768416p pd=3.2364u  as=0.58035p  ps=2.72u   
m05 w4  w2 vdd vdd p w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.382453p ps=1.61081u
m06 vss i2 w2  vss n w=0.54u l=0.13u ad=0.167188p pd=1.23677u as=0.1719p   ps=1.35667u
m07 w2  i1 vss vss n w=0.54u l=0.13u ad=0.1719p   pd=1.35667u as=0.167188p ps=1.23677u
m08 vss i0 w2  vss n w=0.54u l=0.13u ad=0.167188p pd=1.23677u as=0.1719p   ps=1.35667u
m09 nq  w4 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.337473p ps=2.49645u
m10 vss w4 nq  vss n w=1.09u l=0.13u ad=0.337473p pd=2.49645u as=0.28885p  ps=1.62u   
m11 w4  w2 vss vss n w=0.54u l=0.13u ad=0.2295p   pd=1.93u    as=0.167188p ps=1.23677u
C0  vdd w2  0.247f
C1  vdd w1  0.011f
C2  i1  i0  0.224f
C3  i2  w2  0.048f
C4  vdd w3  0.011f
C5  i1  w2  0.028f
C6  vdd nq  0.019f
C7  i0  w4  0.052f
C8  i1  w1  0.012f
C9  i0  w2  0.127f
C10 i1  w3  0.012f
C11 w4  w2  0.146f
C12 vdd i2  0.010f
C13 w2  w1  0.008f
C14 vdd i1  0.010f
C15 w4  nq  0.030f
C16 w2  w3  0.008f
C17 vdd i0  0.030f
C18 w2  nq  0.175f
C19 vdd w4  0.020f
C20 i2  i1  0.257f
C21 nq  vss 0.128f
C22 w3  vss 0.011f
C23 w1  vss 0.011f
C24 w2  vss 0.343f
C25 w4  vss 0.275f
C26 i0  vss 0.137f
C27 i1  vss 0.119f
C28 i2  vss 0.126f
.ends
