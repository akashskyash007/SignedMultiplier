* Spice description of mx3_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:10:33
* ssxlib 0.13um values
.subckt mx3_x2 cmd0 cmd1 i0 i1 i2 q vdd vss
Mtr_00001 vss   cmd1  sig8  vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
Mtr_00002 sig11 cmd0  vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
Mtr_00003 sig1  i1    sig7  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00004 sig7  cmd1  sig6  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00005 sig6  sig8  sig5  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00006 sig5  i2    sig1  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00007 vss   cmd0  sig1  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00008 sig10 sig11 vss   vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00009 sig6  i0    sig10 vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
Mtr_00010 vss   sig6  q     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00011 sig18 sig8  sig6  vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00012 vdd   sig11 sig16 vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00013 sig19 cmd0  vdd   vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00014 sig6  i0    sig19 vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00015 sig16 i1    sig18 vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00016 sig17 i2    sig16 vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00017 sig6  cmd1  sig17 vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00018 q     sig6  vdd   vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00019 sig8  cmd1  vdd   vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
Mtr_00020 vdd   cmd0  sig11 vdd p  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C12 cmd0  vss   1.341f
C3  cmd1  vss   1.550f
C14 i0    vss   0.966f
C9  i1    vss   0.655f
C4  i2    vss   0.545f
C13 q     vss   0.865f
C11 sig11 vss   1.096f
C16 sig16 vss   0.276f
C1  sig1  vss   0.276f
C6  sig6  vss   1.384f
C8  sig8  vss   0.895f
.ends
