.subckt oan21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from oan21_x1.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.1u  l=0.13u ad=0.3883p   pd=2.32667u as=0.41855p  ps=3.06u   
m01 zn  b  vdd vdd p w=0.77u l=0.13u ad=0.20405p  pd=1.372u   as=0.27181p  ps=1.62867u
m02 w1  a2 zn  vdd p w=1.43u l=0.13u ad=0.22165p  pd=1.74u    as=0.37895p  ps=2.548u  
m03 vdd a1 w1  vdd p w=1.43u l=0.13u ad=0.50479p  pd=3.02467u as=0.22165p  ps=1.74u   
m04 z   zn vss vss n w=0.55u l=0.13u ad=0.2002p   pd=1.96u    as=0.208029p ps=1.69706u
m05 n2  b  zn  vss n w=0.66u l=0.13u ad=0.19305p  pd=1.52u    as=0.22935p  ps=2.18u   
m06 vss a2 n2  vss n w=0.66u l=0.13u ad=0.249635p pd=2.03647u as=0.19305p  ps=1.52u   
m07 n2  a1 vss vss n w=0.66u l=0.13u ad=0.19305p  pd=1.52u    as=0.249635p ps=2.03647u
C0  w2  z   0.009f
C1  zn  w3  0.026f
C2  b   n2  0.053f
C3  vdd zn  0.021f
C4  w2  w4  0.166f
C5  w4  w5  0.166f
C6  w2  b   0.011f
C7  z   w3  0.030f
C8  vdd z   0.008f
C9  a2  a1  0.205f
C10 w4  w3  0.166f
C11 w4  vdd 0.051f
C12 w1  w5  0.005f
C13 a2  zn  0.016f
C14 w1  w3  0.001f
C15 a1  zn  0.009f
C16 w4  a2  0.013f
C17 a2  b   0.137f
C18 w4  a1  0.018f
C19 vdd w5  0.020f
C20 a2  w1  0.013f
C21 zn  z   0.136f
C22 a1  b   0.002f
C23 w4  zn  0.031f
C24 vdd w3  0.009f
C25 a2  n2  0.007f
C26 a1  w1  0.012f
C27 zn  b   0.151f
C28 w4  z   0.013f
C29 w2  a2  0.029f
C30 a2  w5  0.002f
C31 a1  n2  0.007f
C32 w4  b   0.018f
C33 a2  w3  0.011f
C34 a1  w5  0.002f
C35 vdd a2  0.002f
C36 w4  w1  0.006f
C37 w2  zn  0.019f
C38 a1  w3  0.011f
C39 zn  w5  0.006f
C40 vdd a1  0.053f
C41 w4  n2  0.036f
C42 w4  vss 1.007f
C43 w2  vss 0.173f
C44 w3  vss 0.163f
C45 w5  vss 0.178f
C46 n2  vss 0.088f
C47 b   vss 0.104f
C48 z   vss 0.040f
C49 zn  vss 0.116f
C50 a1  vss 0.077f
C51 a2  vss 0.096f
.ends
