.subckt nd2v4x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v4x2.ext -        technology: scmos
m00 z   b vdd vdd p w=0.88u  l=0.13u ad=0.1848p    pd=1.3u  as=0.2816p    ps=1.96u
m01 vdd b z   vdd p w=0.88u  l=0.13u ad=0.2816p    pd=1.96u as=0.1848p    ps=1.3u 
m02 z   a vdd vdd p w=0.88u  l=0.13u ad=0.1848p    pd=1.3u  as=0.2816p    ps=1.96u
m03 vdd a z   vdd p w=0.88u  l=0.13u ad=0.2816p    pd=1.96u as=0.1848p    ps=1.3u 
m04 w1  b z   vss n w=0.715u l=0.13u ad=0.0911625p pd=0.97u as=0.268125p  ps=2.18u
m05 vss a w1  vss n w=0.715u l=0.13u ad=0.30745p   pd=2.29u as=0.0911625p ps=0.97u
C0 b   a   0.083f
C1 b   z   0.050f
C2 a   z   0.015f
C3 vdd b   0.003f
C4 vdd a   0.007f
C5 vdd z   0.064f
C6 w1  vss 0.006f
C7 z   vss 0.093f
C8 a   vss 0.151f
C9 b   vss 0.180f
.ends
