* Spice description of vfeed4
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:33
* vsxlib 0.13um values
.subckt vfeed4 vdd vss
.ends
