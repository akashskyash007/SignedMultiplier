.subckt an4v0x2 a b c d vdd vss z
*01-JAN-08 SPICE3       file   created      from an4v0x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.417805p pd=2.76208u as=0.48675p  ps=3.83u   
m01 zn  d  vdd vdd p w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.253667p ps=1.67698u
m02 vdd c  zn  vdd p w=0.935u l=0.13u ad=0.253667p pd=1.67698u as=0.19635p  ps=1.355u  
m03 zn  b  vdd vdd p w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.253667p ps=1.67698u
m04 vdd a  zn  vdd p w=0.935u l=0.13u ad=0.253667p pd=1.67698u as=0.19635p  ps=1.355u  
m05 vss zn z   vss n w=0.77u  l=0.13u ad=0.323627p pd=2.38412u as=0.24035p  ps=2.29u   
m06 w1  d  zn  vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.3278p   ps=2.95u   
m07 w2  c  w1  vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.14025p  ps=1.355u  
m08 w3  b  w2  vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.14025p  ps=1.355u  
m09 vss a  w3  vss n w=1.1u   l=0.13u ad=0.462324p pd=3.40588u as=0.14025p  ps=1.355u  
C0  d  b   0.044f
C1  d  a   0.047f
C2  zn z   0.139f
C3  c  b   0.165f
C4  d  z   0.006f
C5  zn vdd 0.175f
C6  c  a   0.028f
C7  c  z   0.006f
C8  d  vdd 0.007f
C9  b  a   0.182f
C10 c  vdd 0.021f
C11 d  w1  0.009f
C12 b  vdd 0.007f
C13 a  vdd 0.007f
C14 z  vdd 0.034f
C15 w3 a   0.016f
C16 zn d   0.111f
C17 w2 d   0.009f
C18 zn c   0.085f
C19 zn b   0.034f
C20 d  c   0.219f
C21 w3 vss 0.008f
C22 w2 vss 0.011f
C23 w1 vss 0.011f
C25 z  vss 0.237f
C26 a  vss 0.202f
C27 b  vss 0.110f
C28 c  vss 0.112f
C29 d  vss 0.147f
C30 zn vss 0.150f
.ends
