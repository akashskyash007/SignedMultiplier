* Spice description of cgi2v0x05
* Spice driver version 134999461
* Date  1/01/2008 at 16:42:53
* wsclib 0.13um values
.subckt cgi2v0x05 a b c vdd vss z
M01 vdd   a     n1    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 06    a     vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M03 vss   a     n3    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M04 n4    a     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 vdd   b     n1    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M06 z     b     06    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M07 vss   b     n3    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M08 z     b     n4    vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M09 n1    c     z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M10 n3    c     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C4  a     vss   0.874f
C6  b     vss   1.136f
C7  c     vss   0.340f
C9  n1    vss   0.368f
C2  n3    vss   0.280f
C5  z     vss   0.666f
.ends
