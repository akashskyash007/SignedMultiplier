.subckt no4_x4 i0 i1 i2 i3 nq vdd vss
*05-JAN-08 SPICE3       file   created      from no4_x4.ext -        technology: scmos
m00 w1  i1 w2  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=1.18608p  ps=5.59u   
m01 w3  i0 w1  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.32395p  ps=2.4u    
m02 w4  i2 w3  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.32395p  ps=2.4u    
m03 vdd i3 w4  vdd p w=2.09u  l=0.13u ad=0.86151p  pd=3.23559u as=0.32395p  ps=2.4u    
m04 nq  w5 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.884182p ps=3.32074u
m05 vdd w5 nq  vdd p w=2.145u l=0.13u ad=0.884182p pd=3.32074u as=0.568425p ps=2.675u  
m06 w5  w2 vdd vdd p w=1.1u   l=0.13u ad=0.473p    pd=3.06u    as=0.453427p ps=1.70294u
m07 w2  i1 vss vss n w=0.55u  l=0.13u ad=0.148019p pd=1.1075u  as=0.231688p ps=1.43409u
m08 vss i0 w2  vss n w=0.55u  l=0.13u ad=0.231688p pd=1.43409u as=0.148019p ps=1.1075u 
m09 w2  i2 vss vss n w=0.55u  l=0.13u ad=0.148019p pd=1.1075u  as=0.231688p ps=1.43409u
m10 vss i3 w2  vss n w=0.55u  l=0.13u ad=0.231688p pd=1.43409u as=0.148019p ps=1.1075u 
m11 nq  w5 vss vss n w=1.045u l=0.13u ad=0.349525p pd=2.015u   as=0.440206p ps=2.72477u
m12 vss w5 nq  vss n w=1.045u l=0.13u ad=0.440206p pd=2.72477u as=0.349525p ps=2.015u  
m13 w5  w2 vss vss n w=0.55u  l=0.13u ad=0.2365p   pd=1.96u    as=0.231688p ps=1.43409u
C0  i2  w2  0.019f
C1  i3  w5  0.006f
C2  i3  w2  0.019f
C3  i0  w3  0.031f
C4  vdd i1  0.023f
C5  nq  vdd 0.080f
C6  w5  w2  0.210f
C7  vdd i0  0.023f
C8  i2  w4  0.052f
C9  vdd i2  0.023f
C10 vdd i3  0.075f
C11 i1  i0  0.267f
C12 vdd w5  0.051f
C13 i1  i2  0.002f
C14 vdd w2  0.033f
C15 i0  i2  0.275f
C16 vdd w1  0.010f
C17 nq  w5  0.020f
C18 i1  w2  0.215f
C19 vdd w3  0.010f
C20 i2  i3  0.281f
C21 nq  w2  0.095f
C22 i0  w2  0.019f
C23 i1  w1  0.019f
C24 vdd w4  0.010f
C25 nq  vss 0.104f
C26 w4  vss 0.006f
C27 w3  vss 0.009f
C28 w1  vss 0.011f
C29 w2  vss 0.549f
C30 w5  vss 0.328f
C31 i3  vss 0.147f
C32 i2  vss 0.139f
C33 i0  vss 0.149f
C34 i1  vss 0.146f
.ends
