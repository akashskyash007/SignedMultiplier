* Spice description of no2_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:18:19
* sxlib 0.13um values
.subckt no2_x1 i0 i1 nq vdd vss
Mtr_00001 nq    i0    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 vss   i1    nq    vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 sig3  i1    nq    vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00004 vdd   i0    sig3  vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C6  i0    vss   1.009f
C5  i1    vss   0.882f
C1  nq    vss   0.852f
.ends
