.subckt nd2v4x6 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v4x6.ext -        technology: scmos
m00 z   a vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.91u    as=0.37895p  ps=2.44429u
m01 vdd b z   vdd p w=1.43u  l=0.13u ad=0.37895p  pd=2.44429u as=0.3003p   ps=1.91u   
m02 z   b vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.91u    as=0.37895p  ps=2.44429u
m03 vdd a z   vdd p w=1.43u  l=0.13u ad=0.37895p  pd=2.44429u as=0.3003p   ps=1.91u   
m04 z   a vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.91u    as=0.37895p  ps=2.44429u
m05 vdd b z   vdd p w=1.43u  l=0.13u ad=0.37895p  pd=2.44429u as=0.3003p   ps=1.91u   
m06 z   b vdd vdd p w=0.715u l=0.13u ad=0.15015p  pd=0.955u   as=0.189475p ps=1.22214u
m07 vdd a z   vdd p w=0.715u l=0.13u ad=0.189475p pd=1.22214u as=0.15015p  ps=0.955u  
m08 w1  a vss vss n w=1.045u l=0.13u ad=0.133238p pd=1.3u     as=0.591525p ps=3.5u    
m09 z   b w1  vss n w=1.045u l=0.13u ad=0.21945p  pd=1.465u   as=0.133238p ps=1.3u    
m10 w2  b z   vss n w=1.045u l=0.13u ad=0.133238p pd=1.3u     as=0.21945p  ps=1.465u  
m11 vss a w2  vss n w=1.045u l=0.13u ad=0.591525p pd=3.5u     as=0.133238p ps=1.3u    
C0  vdd a   0.021f
C1  vdd b   0.033f
C2  vdd z   0.293f
C3  a   b   0.518f
C4  a   z   0.185f
C5  a   w1  0.006f
C6  b   z   0.142f
C7  a   w2  0.006f
C8  z   w1  0.009f
C9  w2  vss 0.010f
C10 w1  vss 0.008f
C11 z   vss 0.384f
C12 b   vss 0.265f
C13 a   vss 0.343f
.ends
