.subckt iv1v0x2 a vdd vss z
*10-JAN-08 SPICE3       file   created      from iv1v0x2.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 z   a   vdd vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 vss vdd w2  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m03 z   a   vss vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0 a   z   0.167f
C1 vdd a   0.096f
C2 vdd z   0.073f
C3 w2  vss 0.014f
C4 z   vss 0.147f
C5 w1  vss 0.019f
C6 a   vss 0.150f
.ends
