* Spice description of tie_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:41:44
* ssxlib 0.13um values
.subckt tie_x0 vdd vss
.ends
