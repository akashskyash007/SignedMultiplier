.subckt xaoi21_x05 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from xaoi21_x05.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.1u   l=0.13u ad=0.355025p pd=2.015u   as=0.33385p  ps=2.10667u
m01 an  a2 vdd vdd p w=1.1u   l=0.13u ad=0.33385p  pd=2.10667u as=0.355025p ps=2.015u  
m02 z   b  an  vdd p w=1.1u   l=0.13u ad=0.336875p pd=2.29u    as=0.33385p  ps=2.10667u
m03 w1  bn z   vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u    as=0.336875p ps=2.29u   
m04 vdd an w1  vdd p w=1.1u   l=0.13u ad=0.355025p pd=2.015u   as=0.1705p   ps=1.41u   
m05 bn  b  vdd vdd p w=1.1u   l=0.13u ad=0.41855p  pd=3.06u    as=0.355025p ps=2.015u  
m06 w2  a1 vss vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.4411p   ps=3.05714u
m07 an  a2 w2  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.19u    as=0.1023p   ps=0.97u   
m08 z   bn an  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.36u    as=0.1749p   ps=1.19u   
m09 bn  an z   vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u   as=0.131175p ps=1.02u   
m10 vss b  bn  vss n w=0.495u l=0.13u ad=0.330825p pd=2.29286u as=0.131175p ps=1.025u  
C0  a1  w2  0.005f
C1  vdd b   0.144f
C2  bn  an  0.193f
C3  vdd a2  0.014f
C4  bn  b   0.119f
C5  bn  a1  0.009f
C6  an  b   0.207f
C7  bn  a2  0.036f
C8  an  a1  0.128f
C9  bn  z   0.119f
C10 an  a2  0.086f
C11 an  z   0.065f
C12 b   a2  0.032f
C13 an  w1  0.007f
C14 b   z   0.010f
C15 a1  a2  0.163f
C16 an  w2  0.010f
C17 a1  z   0.039f
C18 b   w1  0.012f
C19 vdd bn  0.015f
C20 a2  z   0.067f
C21 vdd an  0.036f
C22 z   vss 0.062f
C23 a2  vss 0.081f
C24 a1  vss 0.106f
C25 b   vss 0.126f
C26 an  vss 0.247f
C27 bn  vss 0.162f
.ends
