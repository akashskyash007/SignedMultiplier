.subckt nr2av0x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2av0x1.ext -        technology: scmos
m00 w1  b  z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.48675p  ps=3.83u   
m01 vdd an w1  vdd p w=1.54u l=0.13u ad=0.5852p   pd=2.77455u as=0.19635p  ps=1.795u  
m02 an  a  vdd vdd p w=0.88u l=0.13u ad=0.31185p  pd=2.51u    as=0.3344p   ps=1.58545u
m03 an  a  vss vss n w=0.44u l=0.13u ad=0.1529p   pd=1.63u    as=0.215417p ps=1.77667u
m04 z   b  vss vss n w=0.44u l=0.13u ad=0.0924p   pd=0.86u    as=0.215417p ps=1.77667u
m05 vss an z   vss n w=0.44u l=0.13u ad=0.215417p pd=1.77667u as=0.0924p   ps=0.86u   
C0  z   a   0.007f
C1  vdd b   0.026f
C2  vdd an  0.012f
C3  vdd z   0.029f
C4  vdd w1  0.004f
C5  b   an  0.137f
C6  vdd a   0.021f
C7  b   z   0.102f
C8  an  z   0.028f
C9  b   w1  0.014f
C10 b   a   0.054f
C11 an  a   0.139f
C12 a   vss 0.110f
C13 w1  vss 0.009f
C14 z   vss 0.289f
C15 an  vss 0.140f
C16 b   vss 0.096f
.ends
