.subckt rowend_x0 vdd vss
*04-JAN-08 SPICE3       file   created      from rowend_x0.ext -        technology: scmos
.ends
