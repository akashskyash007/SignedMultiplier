* Spice description of iv1v1x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:44:44
* vsclib 0.13um values
.subckt iv1v1x2 a vdd vss z
M01 vdd   a     z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M02 vss   a     z     vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C3  a     vss   0.527f
C2  z     vss   0.625f
.ends
