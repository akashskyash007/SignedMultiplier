.subckt xaon21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon21_x1.ext -        technology: scmos
m00 vdd a1 an  vdd p w=2.09u  l=0.13u ad=0.78375p  pd=3.53667u as=0.5962p   ps=3.42667u
m01 an  a2 vdd vdd p w=2.09u  l=0.13u ad=0.5962p   pd=3.42667u as=0.78375p  ps=3.53667u
m02 z   bn an  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.5962p   ps=3.42667u
m03 bn  an z   vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.55385p  ps=2.62u   
m04 vdd b  bn  vdd p w=2.09u  l=0.13u ad=0.78375p  pd=3.53667u as=0.55385p  ps=2.62u   
m05 w1  a1 vss vss n w=1.32u  l=0.13u ad=0.2046p   pd=1.63u    as=0.621095p ps=3.30947u
m06 an  a2 w1  vss n w=1.32u  l=0.13u ad=0.3498p   pd=1.85u    as=0.2046p   ps=1.63u   
m07 z   b  an  vss n w=1.32u  l=0.13u ad=0.37158p  pd=2.22u    as=0.3498p   ps=1.85u   
m08 w2  bn z   vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.24772p  ps=1.48u   
m09 vss an w2  vss n w=0.88u  l=0.13u ad=0.414063p pd=2.20632u as=0.1364p   ps=1.19u   
m10 bn  b  vss vss n w=0.935u l=0.13u ad=0.374825p pd=2.73u    as=0.439942p ps=2.34421u
C0  bn  z   0.016f
C1  an  vdd 0.157f
C2  an  z   0.221f
C3  b   vdd 0.029f
C4  b   z   0.065f
C5  an  w2  0.016f
C6  vdd z   0.017f
C7  a1  a2  0.154f
C8  a1  an  0.011f
C9  a2  bn  0.047f
C10 a2  an  0.088f
C11 bn  an  0.285f
C12 a1  vdd 0.010f
C13 a2  b   0.058f
C14 a2  vdd 0.043f
C15 bn  b   0.157f
C16 a1  z   0.016f
C17 bn  vdd 0.132f
C18 an  b   0.062f
C19 a1  w1  0.013f
C20 w2  vss 0.003f
C21 w1  vss 0.003f
C22 z   vss 0.025f
C24 b   vss 0.229f
C25 an  vss 0.202f
C26 bn  vss 0.152f
C27 a2  vss 0.066f
C28 a1  vss 0.078f
.ends
