.subckt oai21v0x1 a1 a2 b vdd vss z
*10-JAN-08 SPICE3       file   created      from oai21v0x1.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.54u l=0.13u ad=0.537167p pd=3.09667u as=0.5775p   ps=3.83u   
m01 w2  a1  vdd vdd p w=1.54u l=0.13u ad=0.5775p   pd=3.83u    as=0.537167p ps=3.09667u
m02 z   a2  w2  vdd p w=1.54u l=0.13u ad=0.517p    pd=2.73u    as=0.5775p   ps=3.83u   
m03 vdd b   z   vdd p w=1.54u l=0.13u ad=0.537167p pd=3.09667u as=0.517p    ps=2.73u   
m04 vss vdd w3  vss n w=1.1u  l=0.13u ad=0.404433p pd=2.51u    as=0.4125p   ps=2.95u   
m05 w4  a1  vss vss n w=1.1u  l=0.13u ad=0.404433p pd=2.51u    as=0.404433p ps=2.51u   
m06 w4  a2  vss vss n w=1.1u  l=0.13u ad=0.404433p pd=2.51u    as=0.404433p ps=2.51u   
m07 z   b   w4  vss n w=1.1u  l=0.13u ad=0.4125p   pd=2.95u    as=0.404433p ps=2.51u   
C0  vdd z   0.010f
C1  vdd b   0.048f
C2  a1  a2  0.050f
C3  vdd w2  0.017f
C4  a2  z   0.091f
C5  a2  b   0.089f
C6  z   b   0.142f
C7  a1  w2  0.016f
C8  a2  w2  0.016f
C9  z   w2  0.004f
C10 a1  w4  0.006f
C11 a2  w4  0.015f
C12 vdd a1  0.096f
C13 z   w4  0.078f
C14 vdd a2  0.007f
C15 w4  vss 0.151f
C16 w3  vss 0.014f
C17 w2  vss 0.053f
C18 w1  vss 0.019f
C19 b   vss 0.148f
C20 z   vss 0.080f
C21 a2  vss 0.178f
C22 a1  vss 0.155f
.ends
