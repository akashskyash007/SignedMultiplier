.subckt na3_x4 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from na3_x4.ext -        technology: scmos
m00 vdd i0 w1  vdd p w=1.09u l=0.13u ad=0.303392p pd=1.89815u as=0.346983p ps=2.09u   
m01 w1  i2 vdd vdd p w=1.09u l=0.13u ad=0.346983p pd=2.09u    as=0.303392p ps=1.89815u
m02 vdd i1 w1  vdd p w=1.09u l=0.13u ad=0.303392p pd=1.89815u as=0.346983p ps=2.09u   
m03 nq  w2 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.609567p ps=3.81371u
m04 vdd w2 nq  vdd p w=2.19u l=0.13u ad=0.609567p pd=3.81371u as=0.58035p  ps=2.72u   
m05 w2  w1 vdd vdd p w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.303392p ps=1.89815u
m06 w3  i0 w1  vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.46325p  ps=3.03u   
m07 w4  i2 w3  vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.16895p  ps=1.4u    
m08 vss i1 w4  vss n w=1.09u l=0.13u ad=0.415988p pd=2.2315u  as=0.16895p  ps=1.4u    
m09 nq  w2 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.415988p ps=2.2315u 
m10 vss w2 nq  vss n w=1.09u l=0.13u ad=0.415988p pd=2.2315u  as=0.28885p  ps=1.62u   
m11 w2  w1 vss vss n w=0.54u l=0.13u ad=0.2295p   pd=1.93u    as=0.206086p ps=1.10551u
C0  w1  w3  0.008f
C1  i1  w4  0.005f
C2  w1  w4  0.008f
C3  vdd i2  0.019f
C4  w2  i1  0.058f
C5  w2  w1  0.094f
C6  i0  i2  0.222f
C7  w2  nq  0.030f
C8  vdd w1  0.217f
C9  i0  i1  0.005f
C10 i0  w1  0.055f
C11 vdd nq  0.019f
C12 i2  i1  0.216f
C13 i2  w1  0.028f
C14 i1  w1  0.145f
C15 i2  w3  0.009f
C16 w1  nq  0.145f
C17 w2  vdd 0.020f
C18 w4  vss 0.007f
C19 w3  vss 0.006f
C20 nq  vss 0.123f
C21 w1  vss 0.335f
C22 i1  vss 0.138f
C23 i2  vss 0.122f
C24 i0  vss 0.128f
C26 w2  vss 0.277f
.ends
