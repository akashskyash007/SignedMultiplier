* Spice description of oai31v0x1
* Spice driver version 134999461
* Date  1/01/2008 at 16:59:36
* vsclib 0.13um values
.subckt oai31v0x1 a1 a2 a3 b vdd vss z
M01 sig8  a1    vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M02 vdd   a1    05    vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M03 vss   a1    sig1  vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 n2a   a2    sig8  vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M05 05    a2    08    vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M06 vss   a2    sig1  vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M07 z     a3    n2a   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M08 08    a3    z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
M09 sig1  a3    vss   vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M10 vdd   b     z     vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M11 sig1  b     z     vss n  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
C5  a1    vss   1.084f
C6  a2    vss   0.825f
C7  a3    vss   0.515f
C4  b     vss   0.367f
C1  sig1  vss   0.272f
C3  z     vss   0.918f
.ends
