.subckt noa2a2a23_x4 i0 i1 i2 i3 i4 i5 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa2a2a23_x4.ext -        technology: scmos
m00 w1  i5 w2  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.701319p ps=3.83u   
m01 w2  i4 w1  vdd p w=2.09u  l=0.13u ad=0.701319p pd=3.83u    as=0.55385p  ps=2.62u   
m02 w3  i3 w2  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.701319p ps=3.83u   
m03 w2  i2 w3  vdd p w=2.09u  l=0.13u ad=0.701319p pd=3.83u    as=0.55385p  ps=2.62u   
m04 w3  i1 vdd vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.62718p  ps=3.46149u
m05 vdd i0 w3  vdd p w=2.09u  l=0.13u ad=0.62718p  pd=3.46149u as=0.55385p  ps=2.62u   
m06 nq  w4 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.643685p ps=3.55259u
m07 vdd w4 nq  vdd p w=2.145u l=0.13u ad=0.643685p pd=3.55259u as=0.568425p ps=2.675u  
m08 w4  w1 vdd vdd p w=1.1u   l=0.13u ad=0.473p    pd=3.06u    as=0.330095p ps=1.82184u
m09 w5  i5 vss vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.332815p ps=2.11412u
m10 w1  i4 w5  vss n w=0.99u  l=0.13u ad=0.3168p   pd=1.96u    as=0.15345p  ps=1.3u    
m11 w6  i3 w1  vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.3168p   ps=1.96u   
m12 vss i2 w6  vss n w=0.99u  l=0.13u ad=0.332815p pd=2.11412u as=0.15345p  ps=1.3u    
m13 w7  i1 w1  vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.3168p   ps=1.96u   
m14 vss i0 w7  vss n w=0.99u  l=0.13u ad=0.332815p pd=2.11412u as=0.15345p  ps=1.3u    
m15 nq  w4 vss vss n w=1.045u l=0.13u ad=0.349525p pd=2.015u   as=0.351304p ps=2.23157u
m16 vss w4 nq  vss n w=1.045u l=0.13u ad=0.351304p pd=2.23157u as=0.349525p ps=2.015u  
m17 w4  w1 vss vss n w=0.55u  l=0.13u ad=0.2365p   pd=1.96u    as=0.184897p ps=1.17451u
C0  w3  i4  0.009f
C1  w1  i3  0.019f
C2  w2  i2  0.016f
C3  i0  w4  0.094f
C4  w2  w1  0.067f
C5  w1  i2  0.019f
C6  w3  i3  0.024f
C7  w2  w3  0.079f
C8  w1  i1  0.019f
C9  w3  i2  0.019f
C10 i0  vdd 0.010f
C11 vdd i5  0.010f
C12 w3  i1  0.024f
C13 vdd i4  0.010f
C14 w1  nq  0.040f
C15 vdd i3  0.010f
C16 w4  w1  0.159f
C17 w2  vdd 0.179f
C18 vdd i2  0.010f
C19 i5  i4  0.230f
C20 w1  w5  0.010f
C21 w1  vdd 0.017f
C22 vdd i1  0.015f
C23 w4  nq  0.020f
C24 w1  w6  0.010f
C25 w2  i5  0.007f
C26 w3  vdd 0.087f
C27 i4  i3  0.207f
C28 w1  w7  0.010f
C29 i0  w1  0.019f
C30 i0  i1  0.219f
C31 w1  i5  0.163f
C32 w2  i4  0.053f
C33 nq  vdd 0.092f
C34 i0  w3  0.009f
C35 w4  vdd 0.032f
C36 w1  i4  0.030f
C37 w2  i3  0.007f
C38 i3  i2  0.226f
C39 w7  vss 0.014f
C40 w6  vss 0.015f
C41 w5  vss 0.015f
C42 nq  vss 0.096f
C43 w3  vss 0.060f
C44 w1  vss 0.684f
C45 w2  vss 0.104f
C46 w4  vss 0.291f
C47 i0  vss 0.128f
C48 i1  vss 0.135f
C49 i2  vss 0.140f
C50 i3  vss 0.133f
C51 i4  vss 0.148f
C52 i5  vss 0.142f
.ends
