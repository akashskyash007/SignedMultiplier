.subckt xaon22_x05 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon22_x05.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.1u   l=0.13u ad=0.528963p pd=2.1525u  as=0.33385p  ps=2.10667u
m01 an  a2 vdd vdd p w=1.1u   l=0.13u ad=0.33385p  pd=2.10667u as=0.528963p ps=2.1525u 
m02 z   bn an  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.33385p  ps=2.10667u
m03 bn  an z   vdd p w=1.1u   l=0.13u ad=0.414517p pd=2.25333u as=0.2915p   ps=1.63u   
m04 vdd b1 bn  vdd p w=1.1u   l=0.13u ad=0.528963p pd=2.1525u  as=0.414517p ps=2.25333u
m05 bn  b2 vdd vdd p w=1.1u   l=0.13u ad=0.414517p pd=2.25333u as=0.528963p ps=2.1525u 
m06 w1  a1 vss vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.427981p ps=2.38049u
m07 an  a2 w1  vss n w=0.88u  l=0.13u ad=0.2332p   pd=1.41u    as=0.1364p   ps=1.19u   
m08 w2  b2 an  vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.2332p   ps=1.41u   
m09 z   b1 w2  vss n w=0.88u  l=0.13u ad=0.2332p   pd=1.8048u  as=0.1364p   ps=1.19u   
m10 w3  bn z   vss n w=0.495u l=0.13u ad=0.076725p pd=0.805u   as=0.131175p ps=1.0152u 
m11 vss an w3  vss n w=0.495u l=0.13u ad=0.240739p pd=1.33902u as=0.076725p ps=0.805u  
m12 w4  b1 vss vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.427981p ps=2.38049u
m13 bn  b2 w4  vss n w=0.88u  l=0.13u ad=0.28765p  pd=2.62u    as=0.1364p   ps=1.19u   
C0  an  w2  0.010f
C1  a1  a2  0.121f
C2  vdd an  0.105f
C3  an  w3  0.006f
C4  vdd b1  0.028f
C5  a2  bn  0.045f
C6  a1  an  0.007f
C7  z   w2  0.004f
C8  a2  an  0.070f
C9  b2  w4  0.020f
C10 bn  an  0.295f
C11 a2  b2  0.032f
C12 bn  b1  0.110f
C13 a2  z   0.067f
C14 an  b1  0.011f
C15 bn  b2  0.072f
C16 bn  z   0.032f
C17 an  b2  0.009f
C18 an  z   0.203f
C19 b1  b2  0.288f
C20 vdd a2  0.007f
C21 b1  z   0.011f
C22 vdd bn  0.124f
C23 z   vss 0.027f
C24 b2  vss 0.323f
C25 b1  vss 0.190f
C26 an  vss 0.244f
C27 bn  vss 0.150f
C28 a2  vss 0.103f
C29 a1  vss 0.100f
.ends
