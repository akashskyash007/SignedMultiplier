.subckt noa22_x4 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa22_x4.ext -        technology: scmos
m00 w1  i2 vdd vdd p w=1.09u l=0.13u ad=0.346983p pd=2.09u    as=0.428689p ps=2.42259u
m01 w2  i1 w1  vdd p w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.346983p ps=2.09u   
m02 w1  i0 w2  vdd p w=1.09u l=0.13u ad=0.346983p pd=2.09u    as=0.28885p  ps=1.62u   
m03 vdd w2 w3  vdd p w=1.09u l=0.13u ad=0.428689p pd=2.42259u as=0.46325p  ps=3.03u   
m04 nq  w3 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.861311p ps=4.86741u
m05 vdd w3 nq  vdd p w=2.19u l=0.13u ad=0.861311p pd=4.86741u as=0.58035p  ps=2.72u   
m06 w2  i2 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.244961p ps=1.68963u
m07 w4  i1 w2  vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.1431p   ps=1.07u   
m08 vss i0 w4  vss n w=0.54u l=0.13u ad=0.244961p pd=1.68963u as=0.1431p   ps=1.07u   
m09 vss w2 w3  vss n w=0.54u l=0.13u ad=0.244961p pd=1.68963u as=0.2295p   ps=1.93u   
m10 nq  w3 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.494458p ps=3.41055u
m11 vss w3 nq  vss n w=1.09u l=0.13u ad=0.494458p pd=3.41055u as=0.28885p  ps=1.62u   
C0  vdd nq  0.084f
C1  i2  w1  0.010f
C2  w3  w2  0.151f
C3  i1  i0  0.201f
C4  i2  w2  0.119f
C5  w3  nq  0.030f
C6  i1  w1  0.005f
C7  i1  w2  0.114f
C8  i0  w1  0.005f
C9  i0  w2  0.014f
C10 vdd w3  0.020f
C11 i1  w4  0.015f
C12 w1  w2  0.094f
C13 vdd i2  0.046f
C14 vdd i1  0.002f
C15 w2  nq  0.033f
C16 vdd i0  0.002f
C17 vdd w1  0.065f
C18 vdd w2  0.028f
C19 i2  i1  0.076f
C20 w4  vss 0.008f
C21 nq  vss 0.132f
C22 w2  vss 0.186f
C23 w1  vss 0.034f
C24 i0  vss 0.158f
C25 i1  vss 0.171f
C26 i2  vss 0.203f
C27 w3  vss 0.279f
.ends
