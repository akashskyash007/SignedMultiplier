.subckt iv1v6x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v6x2.ext -        technology: scmos
m00 vdd a z vdd p w=1.54u l=0.13u ad=0.810425p pd=4.38u as=0.48675p ps=3.83u
m01 vss a z vss n w=0.77u l=0.13u ad=0.564025p pd=3.5u  as=0.28875p ps=2.29u
C0 vdd a   0.040f
C1 vdd z   0.051f
C2 a   z   0.118f
C3 z   vss 0.232f
C4 a   vss 0.168f
.ends
