.subckt xaoi21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from xaoi21_x1.ext -        technology: scmos
m00 an  a1 vdd vdd p w=2.09u  l=0.13u ad=0.5962p   pd=3.42667u as=0.653675p ps=3.83u   
m01 vdd a2 an  vdd p w=2.09u  l=0.13u ad=0.653675p pd=3.83u    as=0.5962p   ps=3.42667u
m02 z   b  an  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.5962p   ps=3.42667u
m03 w1  bn z   vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.55385p  ps=2.62u   
m04 vdd an w1  vdd p w=2.09u  l=0.13u ad=0.653675p pd=3.83u    as=0.32395p  ps=2.4u    
m05 bn  b  vdd vdd p w=2.09u  l=0.13u ad=0.6809p   pd=5.04u    as=0.653675p ps=3.83u   
m06 w2  a1 vss vss n w=1.32u  l=0.13u ad=0.2046p   pd=1.63u    as=0.652595p ps=3.90439u
m07 an  a2 w2  vss n w=1.32u  l=0.13u ad=0.3498p   pd=1.85u    as=0.2046p   ps=1.63u   
m08 z   bn an  vss n w=1.32u  l=0.13u ad=0.3498p   pd=2.16585u as=0.3498p   ps=1.85u   
m09 bn  an z   vss n w=0.935u l=0.13u ad=0.247775p pd=1.465u   as=0.247775p ps=1.53415u
m10 vss b  bn  vss n w=0.935u l=0.13u ad=0.462255p pd=2.76561u as=0.247775p ps=1.465u  
C0  b   z   0.022f
C1  vdd bn  0.018f
C2  a1  w2  0.008f
C3  b   w1  0.010f
C4  vdd z   0.015f
C5  an  bn  0.265f
C6  an  z   0.185f
C7  vdd w1  0.009f
C8  bn  z   0.020f
C9  an  w1  0.020f
C10 a1  a2  0.202f
C11 an  w2  0.010f
C12 a1  vdd 0.010f
C13 a2  b   0.005f
C14 a1  an  0.132f
C15 a2  vdd 0.022f
C16 b   vdd 0.198f
C17 a1  bn  0.009f
C18 a2  an  0.090f
C19 a2  bn  0.041f
C20 b   an  0.266f
C21 a1  z   0.016f
C22 a2  z   0.012f
C23 vdd an  0.108f
C24 b   bn  0.192f
C25 w2  vss 0.009f
C26 z   vss 0.071f
C27 bn  vss 0.214f
C28 an  vss 0.268f
C30 b   vss 0.160f
C31 a2  vss 0.092f
C32 a1  vss 0.108f
.ends
