* Spice description of iv1v0x4
* Spice driver version 134999461
* Date 10/01/2008 at 16:57:17
* vgalib 0.13um values
.subckt iv1v0x4 a vdd vss z
Mtr_00001 z     a     vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 vss   a     z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 vdd   a     z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00004 z     a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C3  a     vss   1.590f
C2  z     vss   0.581f
.ends
