* Spice description of vfeed1
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:06
* vxlib 0.13um values
.subckt vfeed1 vdd vss
.ends
