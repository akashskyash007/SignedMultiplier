* Spice description of nd2abv0x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:48:47
* wsclib 0.13um values
.subckt nd2abv0x2 a b vdd vss z
M01 sig5  a     vdd   vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M02 sig5  a     vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M03 vdd   b     bn    vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M04 vss   b     bn    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M05 vdd   sig5  z     vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M06 vss   sig5  08    vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M07 z     bn    vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M08 08    bn    z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C7  a     vss   0.490f
C3  bn    vss   0.651f
C4  b     vss   0.557f
C5  sig5  vss   0.587f
C2  z     vss   0.451f
.ends
