.subckt iv1v0x6 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v0x6.ext -        technology: scmos
m00 vdd a z   vdd p w=1.485u l=0.13u ad=0.393525p pd=2.51u  as=0.365292p ps=2.51u 
m01 z   a vdd vdd p w=1.485u l=0.13u ad=0.365292p pd=2.51u  as=0.393525p ps=2.51u 
m02 vdd a z   vdd p w=1.485u l=0.13u ad=0.393525p pd=2.51u  as=0.365292p ps=2.51u 
m03 z   a vss vss n w=1.1u   l=0.13u ad=0.231p    pd=1.52u  as=0.421575p ps=3.005u
m04 vss a z   vss n w=1.1u   l=0.13u ad=0.421575p pd=3.005u as=0.231p    ps=1.52u 
C0 z vdd 0.025f
C1 a z   0.076f
C2 a vdd 0.035f
C4 z vss 0.261f
C5 a vss 0.251f
.ends
