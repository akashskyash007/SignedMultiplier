* Spice description of nd2v6x4
* Spice driver version 134999461
* Date 10/01/2008 at 16:57:46
* vgalib 0.13um values
.subckt nd2v6x4 a b vdd vss z
Mtr_00001 z     b     sig1  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00002 sig1  b     z     vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00003 sig1  a     vss   vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00004 vss   a     sig1  vss n  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
Mtr_00005 vdd   b     z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00006 z     b     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00007 vdd   a     z     vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
Mtr_00008 z     a     vdd   vdd p  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C3  a     vss   1.460f
C5  b     vss   1.528f
C1  sig1  vss   0.275f
C4  z     vss   1.060f
.ends
