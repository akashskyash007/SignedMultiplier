.subckt iv1v0x6 a vdd vss z
*10-JAN-08 SPICE3       file   created      from iv1v0x6.ext -        technology: scmos
m00 z   a   vdd vdd p w=1.43u l=0.13u ad=0.37895p pd=1.96u as=0.53625p ps=3.61u
m01 vdd a   z   vdd p w=1.43u l=0.13u ad=0.53625p pd=3.61u as=0.37895p ps=1.96u
m02 z   a   vdd vdd p w=1.43u l=0.13u ad=0.37895p pd=1.96u as=0.53625p ps=3.61u
m03 w1  vdd z   vdd p w=1.43u l=0.13u ad=0.53625p pd=3.61u as=0.37895p ps=1.96u
m04 z   a   vss vss n w=0.99u l=0.13u ad=0.26235p pd=1.52u as=0.37125p ps=2.73u
m05 vss a   z   vss n w=0.99u l=0.13u ad=0.37125p pd=2.73u as=0.26235p ps=1.52u
m06 z   a   vss vss n w=0.99u l=0.13u ad=0.26235p pd=1.52u as=0.37125p ps=2.73u
m07 w2  vss z   vss n w=0.99u l=0.13u ad=0.37125p pd=2.73u as=0.26235p ps=1.52u
C0 vdd a   0.106f
C1 vdd z   0.091f
C2 a   z   0.159f
C3 w2  vss 0.011f
C4 w1  vss 0.014f
C5 z   vss 0.261f
C6 a   vss 0.697f
.ends
