.subckt ha2_x2 a b co so vdd vss
*04-JAN-08 SPICE3       file   created      from ha2_x2.ext -        technology: scmos
m00 vdd son so  vdd p w=2.09u  l=0.13u ad=0.637245p pd=2.96922u as=0.6809p   ps=5.04u   
m01 son con vdd vdd p w=0.99u  l=0.13u ad=0.26235p  pd=1.66154u as=0.301853p ps=1.40647u
m02 w1  b   son vdd p w=1.87u  l=0.13u ad=0.28985p  pd=2.18u    as=0.49555p  ps=3.13846u
m03 vdd a   w1  vdd p w=1.87u  l=0.13u ad=0.570167p pd=2.65667u as=0.28985p  ps=2.18u   
m04 con a   vdd vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.637245p ps=2.96922u
m05 vdd b   con vdd p w=2.09u  l=0.13u ad=0.637245p pd=2.96922u as=0.55385p  ps=2.62u   
m06 co  con vdd vdd p w=2.09u  l=0.13u ad=0.6809p   pd=5.04u    as=0.637245p ps=2.96922u
m07 vss son so  vss n w=1.045u l=0.13u ad=0.326286p pd=2.02294u as=0.403975p ps=2.95u   
m08 n2  con vss vss n w=0.825u l=0.13u ad=0.236775p pd=1.74u    as=0.257594p ps=1.59706u
m09 son b   n2  vss n w=0.825u l=0.13u ad=0.232238p pd=1.52u    as=0.236775p ps=1.74u   
m10 n2  a   son vss n w=0.825u l=0.13u ad=0.236775p pd=1.74u    as=0.232238p ps=1.52u   
m11 w2  a   con vss n w=1.76u  l=0.13u ad=0.2728p   pd=2.07u    as=0.52085p  ps=4.38u   
m12 vss b   w2  vss n w=1.76u  l=0.13u ad=0.549534p pd=3.40706u as=0.2728p   ps=2.07u   
m13 co  con vss vss n w=1.045u l=0.13u ad=0.403975p pd=2.95u    as=0.326286p ps=2.02294u
C0  w3  son 0.039f
C1  w4  so  0.014f
C2  w5  vdd 0.040f
C3  n2  a   0.024f
C4  b   con 0.347f
C5  w6  son 0.034f
C6  w3  so  0.009f
C7  w4  vdd 0.013f
C8  w5  b   0.005f
C9  a   con 0.033f
C10 w1  w6  0.004f
C11 co  vdd 0.009f
C12 w6  so  0.036f
C13 w4  b   0.059f
C14 w5  a   0.005f
C15 w2  con 0.010f
C16 w6  vdd 0.074f
C17 w4  a   0.001f
C18 w3  b   0.019f
C19 w5  con 0.017f
C20 son so  0.043f
C21 w6  b   0.025f
C22 w3  a   0.017f
C23 w4  con 0.022f
C24 son vdd 0.015f
C25 co  con 0.179f
C26 w2  w3  0.001f
C27 n2  w6  0.054f
C28 w1  vdd 0.005f
C29 w6  a   0.027f
C30 w3  con 0.012f
C31 so  vdd 0.009f
C32 son b   0.108f
C33 co  w5  0.004f
C34 w2  w6  0.010f
C35 w6  con 0.065f
C36 w1  b   0.012f
C37 n2  son 0.070f
C38 son a   0.009f
C39 co  w4  0.012f
C40 w5  w6  0.166f
C41 vdd b   0.042f
C42 son con 0.210f
C43 co  w3  0.009f
C44 w4  w6  0.166f
C45 w1  con 0.010f
C46 w5  son 0.006f
C47 so  con 0.049f
C48 vdd a   0.018f
C49 co  w6  0.034f
C50 w3  w6  0.166f
C51 w1  w5  0.005f
C52 w4  son 0.018f
C53 w5  so  0.004f
C54 n2  b   0.007f
C55 vdd con 0.177f
C56 b   a   0.378f
C57 w6  vss 0.907f
C58 w3  vss 0.160f
C59 w4  vss 0.143f
C60 w5  vss 0.152f
C61 w2  vss 0.010f
C62 n2  vss 0.094f
C63 co  vss 0.041f
C64 con vss 0.194f
C65 a   vss 0.158f
C66 b   vss 0.154f
C68 so  vss 0.031f
C69 son vss 0.100f
.ends
