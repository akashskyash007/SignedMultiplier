.subckt iv1v5x6 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v5x6.ext -        technology: scmos
m00 vdd a z   vdd p w=1.54u l=0.13u ad=0.4081p   pd=2.58333u as=0.37785p  ps=2.58333u
m01 z   a vdd vdd p w=1.54u l=0.13u ad=0.37785p  pd=2.58333u as=0.4081p   ps=2.58333u
m02 vdd a z   vdd p w=1.54u l=0.13u ad=0.4081p   pd=2.58333u as=0.37785p  ps=2.58333u
m03 z   a vss vss n w=0.88u l=0.13u ad=0.1848p   pd=1.3u     as=0.325463p ps=2.51u   
m04 vss a z   vss n w=0.88u l=0.13u ad=0.325463p pd=2.51u    as=0.1848p   ps=1.3u    
C0 z vdd 0.027f
C1 a z   0.115f
C2 a vdd 0.021f
C4 z vss 0.221f
C5 a vss 0.205f
.ends
