.subckt nd4v0x2 a b c d vdd vss z
*01-JAN-08 SPICE3       file   created      from nd4v0x2.ext -        technology: scmos
m00 z   a vdd vdd p w=1.375u l=0.13u ad=0.28875p  pd=1.795u  as=0.486888p ps=2.8125u
m01 vdd b z   vdd p w=1.375u l=0.13u ad=0.486888p pd=2.8125u as=0.28875p  ps=1.795u 
m02 z   c vdd vdd p w=1.375u l=0.13u ad=0.28875p  pd=1.795u  as=0.486888p ps=2.8125u
m03 vdd d z   vdd p w=1.375u l=0.13u ad=0.486888p pd=2.8125u as=0.28875p  ps=1.795u 
m04 w1  a vss vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.419788p ps=2.785u 
m05 w2  b w1  vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.105188p ps=1.08u  
m06 w3  c w2  vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.105188p ps=1.08u  
m07 z   d w3  vss n w=0.825u l=0.13u ad=0.17325p  pd=1.245u  as=0.105188p ps=1.08u  
m08 w4  d z   vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.17325p  ps=1.245u 
m09 w5  c w4  vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.105188p ps=1.08u  
m10 w6  b w5  vss n w=0.825u l=0.13u ad=0.105188p pd=1.08u   as=0.105188p ps=1.08u  
m11 vss a w6  vss n w=0.825u l=0.13u ad=0.419788p pd=2.785u  as=0.105188p ps=1.08u  
C0  vdd b   0.107f
C1  w4  a   0.002f
C2  z   w1  0.009f
C3  vdd c   0.022f
C4  z   w2  0.009f
C5  vdd d   0.007f
C6  a   b   0.204f
C7  vdd z   0.194f
C8  a   c   0.081f
C9  w3  a   0.002f
C10 a   d   0.125f
C11 b   c   0.330f
C12 a   z   0.201f
C13 b   d   0.105f
C14 b   z   0.116f
C15 c   d   0.306f
C16 w5  a   0.010f
C17 a   w1  0.002f
C18 c   z   0.020f
C19 w3  z   0.009f
C20 w6  a   0.003f
C21 a   w2  0.002f
C22 d   z   0.013f
C23 vdd a   0.007f
C24 w6  vss 0.009f
C25 w5  vss 0.007f
C26 w4  vss 0.010f
C27 w3  vss 0.008f
C28 w2  vss 0.008f
C29 w1  vss 0.009f
C30 z   vss 0.358f
C31 d   vss 0.164f
C32 c   vss 0.176f
C33 b   vss 0.240f
C34 a   vss 0.225f
.ends
