* Spice description of vfeed7
* Spice driver version 134999461
* Date  1/01/2008 at 17:03:03
* vsclib 0.13um values
.subckt vfeed7 vdd vss
.ends
