.subckt o4_x2 i0 i1 i2 i3 q vdd vss
*05-JAN-08 SPICE3       file   created      from o4_x2.ext -        technology: scmos
m00 w1  i3 w2  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.697p    ps=4.13u   
m01 w3  i1 w1  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.2542p   ps=1.95u   
m02 w4  i0 w3  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.2542p   ps=1.95u   
m03 vdd i2 w4  vdd p w=1.64u l=0.13u ad=0.988047p pd=2.80042u as=0.2542p   ps=1.95u   
m04 q   w2 vdd vdd p w=2.19u l=0.13u ad=0.93075p  pd=5.23u    as=1.3194p   ps=3.73958u
m05 w2  i3 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.208631p ps=1.54357u
m06 vss i1 w2  vss n w=0.54u l=0.13u ad=0.208631p pd=1.54357u as=0.1431p   ps=1.07u   
m07 w2  i0 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.208631p ps=1.54357u
m08 vss i2 w2  vss n w=0.54u l=0.13u ad=0.208631p pd=1.54357u as=0.1431p   ps=1.07u   
m09 q   w2 vss vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.421126p ps=3.11572u
C0  i1  w3  0.012f
C1  w2  q   0.238f
C2  w2  i0  0.028f
C3  i3  i1  0.240f
C4  w2  i2  0.154f
C5  i0  w4  0.020f
C6  i1  i0  0.234f
C7  w2  w1  0.008f
C8  i1  w1  0.012f
C9  i0  i2  0.232f
C10 vdd w2  0.174f
C11 vdd i3  0.002f
C12 vdd i1  0.002f
C13 w2  w3  0.008f
C14 vdd q   0.036f
C15 vdd i0  0.002f
C16 w2  i3  0.034f
C17 w2  w4  0.008f
C18 w2  i1  0.029f
C19 vdd i2  0.036f
C20 q   vss 0.119f
C21 w4  vss 0.011f
C22 w3  vss 0.010f
C23 w1  vss 0.010f
C24 i2  vss 0.134f
C25 i0  vss 0.130f
C26 i1  vss 0.119f
C27 i3  vss 0.127f
C28 w2  vss 0.328f
.ends
