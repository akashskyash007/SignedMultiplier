.subckt xaon22_x05 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon22_x05.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.1u   l=0.13u ad=0.528963p pd=2.1525u  as=0.33385p  ps=2.10667u
m01 an  a2 vdd vdd p w=1.1u   l=0.13u ad=0.33385p  pd=2.10667u as=0.528963p ps=2.1525u 
m02 z   bn an  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.33385p  ps=2.10667u
m03 bn  an z   vdd p w=1.1u   l=0.13u ad=0.414517p pd=2.25333u as=0.2915p   ps=1.63u   
m04 vdd b1 bn  vdd p w=1.1u   l=0.13u ad=0.528963p pd=2.1525u  as=0.414517p ps=2.25333u
m05 bn  b2 vdd vdd p w=1.1u   l=0.13u ad=0.414517p pd=2.25333u as=0.528963p ps=2.1525u 
m06 w1  a1 vss vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.427981p ps=2.38049u
m07 an  a2 w1  vss n w=0.88u  l=0.13u ad=0.2332p   pd=1.41u    as=0.1364p   ps=1.19u   
m08 w2  b2 an  vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.2332p   ps=1.41u   
m09 z   b1 w2  vss n w=0.88u  l=0.13u ad=0.2332p   pd=1.8048u  as=0.1364p   ps=1.19u   
m10 w3  bn z   vss n w=0.495u l=0.13u ad=0.076725p pd=0.805u   as=0.131175p ps=1.0152u 
m11 vss an w3  vss n w=0.495u l=0.13u ad=0.240739p pd=1.33902u as=0.076725p ps=0.805u  
m12 w4  b1 vss vss n w=0.88u  l=0.13u ad=0.1364p   pd=1.19u    as=0.427981p ps=2.38049u
m13 bn  b2 w4  vss n w=0.88u  l=0.13u ad=0.28765p  pd=2.62u    as=0.1364p   ps=1.19u   
C0  a1  an  0.007f
C1  a2  bn  0.045f
C2  b2  w5  0.051f
C3  z   an  0.203f
C4  w2  w5  0.005f
C5  w5  b1  0.023f
C6  a2  an  0.070f
C7  z   w2  0.004f
C8  z   b1  0.011f
C9  b2  a2  0.032f
C10 w3  w5  0.002f
C11 w6  vdd 0.019f
C12 bn  an  0.295f
C13 b2  bn  0.072f
C14 w4  w5  0.001f
C15 w7  vdd 0.001f
C16 bn  b1  0.110f
C17 b2  an  0.009f
C18 w6  w5  0.166f
C19 w6  a1  0.002f
C20 w2  an  0.010f
C21 an  b1  0.011f
C22 z   w6  0.006f
C23 b2  b1  0.288f
C24 w7  w5  0.166f
C25 w5  vdd 0.067f
C26 w7  a1  0.002f
C27 w6  a2  0.002f
C28 w3  an  0.006f
C29 z   w7  0.013f
C30 w8  w5  0.166f
C31 w8  a1  0.030f
C32 w7  a2  0.030f
C33 w6  bn  0.044f
C34 z   w8  0.009f
C35 vdd a2  0.007f
C36 b2  w4  0.020f
C37 w5  a1  0.018f
C38 w8  a2  0.009f
C39 w7  bn  0.020f
C40 w6  an  0.016f
C41 z   w5  0.024f
C42 vdd bn  0.124f
C43 b2  w6  0.001f
C44 w6  b1  0.001f
C45 w5  a2  0.018f
C46 w8  bn  0.010f
C47 w7  an  0.014f
C48 vdd an  0.105f
C49 a1  a2  0.121f
C50 b2  w7  0.002f
C51 z   a2  0.067f
C52 w5  bn  0.039f
C53 w8  an  0.017f
C54 w7  b1  0.032f
C55 vdd b1  0.028f
C56 b2  w8  0.023f
C57 z   bn  0.032f
C58 w1  w5  0.007f
C59 w5  an  0.096f
C60 w8  b1  0.001f
C61 w5  vss 0.934f
C62 w8  vss 0.166f
C63 w7  vss 0.158f
C64 w6  vss 0.152f
C65 z   vss 0.027f
C66 b2  vss 0.323f
C67 b1  vss 0.190f
C68 an  vss 0.244f
C69 bn  vss 0.150f
C70 a2  vss 0.103f
C71 a1  vss 0.100f
.ends
