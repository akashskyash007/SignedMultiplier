.subckt cgi2_x2 a b c vdd vss z
*04-JAN-08 SPICE3       file   created      from cgi2_x2.ext -        technology: scmos
m00 n2  a vdd vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.669854p ps=3.37167u
m01 z   c n2  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.539275p ps=2.565u  
m02 n2  c z   vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.539275p ps=2.565u  
m03 vdd a n2  vdd p w=2.035u l=0.13u ad=0.669854p pd=3.37167u as=0.539275p ps=2.565u  
m04 w1  a vdd vdd p w=2.035u l=0.13u ad=0.315425p pd=2.345u   as=0.669854p ps=3.37167u
m05 z   b w1  vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.315425p ps=2.345u  
m06 w2  b z   vdd p w=2.035u l=0.13u ad=0.315425p pd=2.345u   as=0.539275p ps=2.565u  
m07 vdd a w2  vdd p w=2.035u l=0.13u ad=0.669854p pd=3.37167u as=0.315425p ps=2.345u  
m08 n2  b vdd vdd p w=2.035u l=0.13u ad=0.539275p pd=2.565u   as=0.669854p ps=3.37167u
m09 vdd b n2  vdd p w=2.035u l=0.13u ad=0.669854p pd=3.37167u as=0.539275p ps=2.565u  
m10 n4  a vss vss n w=1.815u l=0.13u ad=0.480975p pd=3.0954u  as=0.893252p ps=4.1844u 
m11 z   c n4  vss n w=0.935u l=0.13u ad=0.247775p pd=1.465u   as=0.247775p ps=1.5946u 
m12 n4  c z   vss n w=0.935u l=0.13u ad=0.247775p pd=1.5946u  as=0.247775p ps=1.465u  
m13 vss b n4  vss n w=1.815u l=0.13u ad=0.893252p pd=4.1844u  as=0.480975p ps=3.0954u 
m14 w3  a vss vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u   as=0.46016p  ps=2.1556u 
m15 z   b w3  vss n w=0.935u l=0.13u ad=0.247775p pd=1.465u   as=0.144925p ps=1.245u  
m16 w4  b z   vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u   as=0.247775p ps=1.465u  
m17 vss a w4  vss n w=0.935u l=0.13u ad=0.46016p  pd=2.1556u  as=0.144925p ps=1.245u  
C0  a   z   0.243f
C1  c   n2  0.026f
C2  b   vdd 0.041f
C3  c   z   0.066f
C4  a   w1  0.010f
C5  b   n2  0.020f
C6  b   z   0.169f
C7  a   w2  0.010f
C8  vdd n2  0.366f
C9  vdd z   0.052f
C10 c   n4  0.043f
C11 n2  z   0.053f
C12 vdd w1  0.010f
C13 n2  w1  0.010f
C14 vdd w2  0.010f
C15 z   w1  0.010f
C16 n2  w2  0.010f
C17 a   c   0.215f
C18 a   b   0.520f
C19 z   n4  0.087f
C20 a   vdd 0.098f
C21 c   b   0.026f
C22 z   w3  0.010f
C23 a   n2  0.265f
C24 c   vdd 0.020f
C25 w4  vss 0.011f
C26 w3  vss 0.009f
C27 n4  vss 0.158f
C28 w2  vss 0.010f
C29 w1  vss 0.008f
C30 z   vss 0.219f
C31 n2  vss 0.139f
C33 b   vss 0.446f
C34 c   vss 0.197f
C35 a   vss 0.384f
.ends
