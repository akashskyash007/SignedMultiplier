.subckt vfeed2 vdd vss
*04-JAN-08 SPICE3       file   created      from vfeed2.ext -        technology: scmos
.ends
