.subckt nr2v0x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2v0x1.ext -        technology: scmos
m00 w1  b z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u as=0.48675p  ps=3.83u 
m01 vdd a w1  vdd p w=1.54u l=0.13u ad=0.7469p   pd=4.05u  as=0.19635p  ps=1.795u
m02 z   b vss vss n w=0.44u l=0.13u ad=0.118113p pd=1.08u  as=0.258775p ps=2.18u 
m03 vss a z   vss n w=0.44u l=0.13u ad=0.258775p pd=2.18u  as=0.118113p ps=1.08u 
C0  b  a   0.137f
C1  b  z   0.057f
C2  b  w1  0.006f
C3  a  z   0.008f
C4  b  vdd 0.011f
C5  a  vdd 0.007f
C6  z  vdd 0.020f
C7  w1 vdd 0.004f
C9  w1 vss 0.010f
C10 z  vss 0.282f
C11 a  vss 0.100f
C12 b  vss 0.084f
.ends
