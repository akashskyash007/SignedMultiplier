.subckt one_x0 q vdd vss
*05-JAN-08 SPICE3       file   created      from one_x0.ext -        technology: scmos
m00 q vss vdd vdd p w=1.09u l=0.13u ad=0.46325p pd=3.03u as=0.58315p ps=3.25u
C0 vdd q   0.057f
C1 q   vss 0.191f
.ends
