.subckt oai21v0x1 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from oai21v0x1.ext -        technology: scmos
m00 z   b  vdd vdd p w=0.77u  l=0.13u ad=0.175128p pd=1.30098u as=0.303211p ps=2.08976u
m01 w1  a2 z   vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.337747p ps=2.50902u
m02 vdd a1 w1  vdd p w=1.485u l=0.13u ad=0.584764p pd=4.03024u as=0.189338p ps=1.74u   
m03 n1  b  z   vss n w=0.66u  l=0.13u ad=0.1628p   pd=1.41u    as=0.2112p   ps=2.07u   
m04 vss a2 n1  vss n w=0.66u  l=0.13u ad=0.1386p   pd=1.08u    as=0.1628p   ps=1.41u   
m05 n1  a1 vss vss n w=0.66u  l=0.13u ad=0.1628p   pd=1.41u    as=0.1386p   ps=1.08u   
C0  a1  n1  0.024f
C1  z   n1  0.016f
C2  vdd b   0.007f
C3  vdd a2  0.007f
C4  vdd a1  0.007f
C5  vdd z   0.095f
C6  b   a2  0.143f
C7  b   a1  0.011f
C8  vdd w1  0.004f
C9  b   z   0.108f
C10 a2  a1  0.181f
C11 a2  z   0.020f
C12 b   n1  0.039f
C13 a2  w1  0.015f
C14 a2  n1  0.006f
C15 n1  vss 0.137f
C16 w1  vss 0.006f
C17 z   vss 0.211f
C18 a1  vss 0.111f
C19 a2  vss 0.104f
C20 b   vss 0.128f
.ends
