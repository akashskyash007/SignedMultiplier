.subckt oan21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from oan21_x1.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.1u  l=0.13u ad=0.3883p   pd=2.32667u as=0.41855p  ps=3.06u   
m01 zn  b  vdd vdd p w=0.77u l=0.13u ad=0.20405p  pd=1.372u   as=0.27181p  ps=1.62867u
m02 w1  a2 zn  vdd p w=1.43u l=0.13u ad=0.22165p  pd=1.74u    as=0.37895p  ps=2.548u  
m03 vdd a1 w1  vdd p w=1.43u l=0.13u ad=0.50479p  pd=3.02467u as=0.22165p  ps=1.74u   
m04 z   zn vss vss n w=0.55u l=0.13u ad=0.2002p   pd=1.96u    as=0.208029p ps=1.69706u
m05 n2  b  zn  vss n w=0.66u l=0.13u ad=0.19305p  pd=1.52u    as=0.22935p  ps=2.18u   
m06 vss a2 n2  vss n w=0.66u l=0.13u ad=0.249635p pd=2.03647u as=0.19305p  ps=1.52u   
m07 n2  a1 vss vss n w=0.66u l=0.13u ad=0.19305p  pd=1.52u    as=0.249635p ps=2.03647u
C0  a2  n2  0.007f
C1  a1  w1  0.012f
C2  zn  b   0.151f
C3  a1  n2  0.007f
C4  vdd a2  0.002f
C5  vdd a1  0.053f
C6  b   n2  0.053f
C7  vdd zn  0.021f
C8  vdd z   0.008f
C9  a2  a1  0.205f
C10 a2  zn  0.016f
C11 a1  zn  0.009f
C12 a2  b   0.137f
C13 a2  w1  0.013f
C14 zn  z   0.136f
C15 a1  b   0.002f
C16 n2  vss 0.124f
C17 w1  vss 0.011f
C18 b   vss 0.134f
C19 z   vss 0.092f
C20 zn  vss 0.198f
C21 a1  vss 0.109f
C22 a2  vss 0.151f
.ends
