.subckt aon21bv0x3 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from aon21bv0x3.ext -        technology: scmos
m00 z   an vdd vdd p w=0.935u l=0.13u ad=0.19635p   pd=1.355u   as=0.269129p  ps=1.80517u
m01 vdd b  z   vdd p w=0.935u l=0.13u ad=0.269129p  pd=1.80517u as=0.19635p   ps=1.355u  
m02 z   b  vdd vdd p w=0.935u l=0.13u ad=0.19635p   pd=1.355u   as=0.269129p  ps=1.80517u
m03 vdd an z   vdd p w=0.935u l=0.13u ad=0.269129p  pd=1.80517u as=0.19635p   ps=1.355u  
m04 an  a1 vdd vdd p w=1.375u l=0.13u ad=0.28875p   pd=1.795u   as=0.395779p  ps=2.65466u
m05 vdd a2 an  vdd p w=1.375u l=0.13u ad=0.395779p  pd=2.65466u as=0.28875p   ps=1.795u  
m06 w1  an vss vss n w=0.605u l=0.13u ad=0.0771375p pd=0.86u    as=0.255297p  ps=1.54917u
m07 z   b  w1  vss n w=0.605u l=0.13u ad=0.13418p   pd=1.06464u as=0.0771375p ps=0.86u   
m08 w2  b  z   vss n w=0.935u l=0.13u ad=0.119213p  pd=1.19u    as=0.20737p   ps=1.64536u
m09 vss an w2  vss n w=0.935u l=0.13u ad=0.394551p  pd=2.39417u as=0.119213p  ps=1.19u   
m10 w3  a1 vss vss n w=1.1u   l=0.13u ad=0.14025p   pd=1.355u   as=0.464177p  ps=2.81667u
m11 an  a2 w3  vss n w=1.1u   l=0.13u ad=0.3278p    pd=2.95u    as=0.14025p   ps=1.355u  
C0  an  w3  0.008f
C1  vdd z   0.083f
C2  a1  w3  0.008f
C3  z   w1  0.005f
C4  an  b   0.286f
C5  an  a1  0.195f
C6  an  a2  0.042f
C7  an  vdd 0.076f
C8  an  z   0.163f
C9  b   vdd 0.011f
C10 a1  a2  0.152f
C11 an  w1  0.005f
C12 b   z   0.085f
C13 a1  vdd 0.009f
C14 an  w2  0.005f
C15 a2  vdd 0.006f
C16 w3  vss 0.010f
C17 w2  vss 0.007f
C18 w1  vss 0.002f
C19 z   vss 0.318f
C21 a2  vss 0.115f
C22 a1  vss 0.100f
C23 b   vss 0.152f
C24 an  vss 0.354f
.ends
