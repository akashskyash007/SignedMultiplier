.subckt powmid_x0 vdd vss
*05-JAN-08 SPICE3       file   created      from powmid_x0.ext -        technology: scmos
.ends
