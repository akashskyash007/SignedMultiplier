.subckt on12_x4 i0 i1 q vdd vss
*05-JAN-08 SPICE3       file   created      from on12_x4.ext -        technology: scmos
m00 vdd i0 w1  vdd p w=1.09u l=0.13u ad=0.382795p pd=2.10028u as=0.46325p  ps=3.03u   
m01 w2  w1 w3  vdd p w=1.64u l=0.13u ad=0.2542p   pd=1.95u    as=0.697p    ps=4.13u   
m02 vdd i1 w2  vdd p w=1.64u l=0.13u ad=0.575949p pd=3.16006u as=0.2542p   ps=1.95u   
m03 q   w3 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.769103p ps=4.21983u
m04 vdd w3 q   vdd p w=2.19u l=0.13u ad=0.769103p pd=4.21983u as=0.58035p  ps=2.72u   
m05 vss i0 w1  vss n w=0.54u l=0.13u ad=0.261673p pd=1.44521u as=0.2295p   ps=1.93u   
m06 w3  w1 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.261673p ps=1.44521u
m07 vss i1 w3  vss n w=0.54u l=0.13u ad=0.261673p pd=1.44521u as=0.1431p   ps=1.07u   
m08 q   w3 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.528191p ps=2.91718u
m09 vss w3 q   vss n w=1.09u l=0.13u ad=0.528191p pd=2.91718u as=0.28885p  ps=1.62u   
C0  w3  w2  0.004f
C1  w3  q   0.007f
C2  i1  q   0.166f
C3  vdd i0  0.030f
C4  vdd w1  0.028f
C5  vdd w3  0.031f
C6  vdd i1  0.064f
C7  i0  w1  0.125f
C8  i0  w3  0.060f
C9  vdd q   0.076f
C10 w1  w3  0.027f
C11 w1  i1  0.089f
C12 w3  i1  0.193f
C13 q   vss 0.137f
C14 w2  vss 0.014f
C15 i1  vss 0.172f
C16 w3  vss 0.302f
C17 w1  vss 0.306f
C18 i0  vss 0.196f
.ends
