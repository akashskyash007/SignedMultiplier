.subckt bf1v2x8 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v2x8.ext -        technology: scmos
m00 z   an vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.85u    as=0.380013p ps=2.43311u
m01 vdd an z   vdd p w=1.43u  l=0.13u ad=0.380013p pd=2.43311u as=0.3003p   ps=1.85u   
m02 z   an vdd vdd p w=1.43u  l=0.13u ad=0.3003p   pd=1.85u    as=0.380013p ps=2.43311u
m03 vdd an z   vdd p w=1.43u  l=0.13u ad=0.380013p pd=2.43311u as=0.3003p   ps=1.85u   
m04 an  a  vdd vdd p w=1.43u  l=0.13u ad=0.3146p   pd=2.18636u as=0.380013p ps=2.43311u
m05 vdd a  an  vdd p w=0.99u  l=0.13u ad=0.263086p pd=1.68446u as=0.2178p   ps=1.51364u
m06 z   an vss vss n w=0.715u l=0.13u ad=0.15015p  pd=1.135u   as=0.196383p ps=1.54419u
m07 vss an z   vss n w=0.715u l=0.13u ad=0.196383p pd=1.54419u as=0.15015p  ps=1.135u  
m08 z   an vss vss n w=0.715u l=0.13u ad=0.15015p  pd=1.135u   as=0.196383p ps=1.54419u
m09 vss an z   vss n w=0.715u l=0.13u ad=0.196383p pd=1.54419u as=0.15015p  ps=1.135u  
m10 an  a  vss vss n w=0.605u l=0.13u ad=0.12705p  pd=1.025u   as=0.166171p ps=1.30662u
m11 vss a  an  vss n w=0.605u l=0.13u ad=0.166171p pd=1.30662u as=0.12705p  ps=1.025u  
C0 vdd z   0.031f
C1 an  a   0.144f
C2 an  z   0.178f
C3 vdd an  0.031f
C4 vdd a   0.026f
C5 z   vss 0.281f
C6 a   vss 0.160f
C7 an  vss 0.329f
.ends
