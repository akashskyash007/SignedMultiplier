.subckt bf1v1x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v1x2.ext -        technology: scmos
m00 vdd an z   vdd p w=1.54u  l=0.13u ad=0.470213p pd=2.576u as=0.48675p  ps=3.83u 
m01 an  a  vdd vdd p w=0.935u l=0.13u ad=0.284075p pd=2.62u  as=0.285487p ps=1.564u
m02 vss an z   vss n w=1.045u l=0.13u ad=0.322905p pd=1.995u as=0.355575p ps=2.84u 
m03 an  a  vss vss n w=0.605u l=0.13u ad=0.196625p pd=1.96u  as=0.186945p ps=1.155u
C0 vdd an  0.039f
C1 vdd z   0.054f
C2 an  z   0.133f
C3 an  a   0.156f
C4 a   vss 0.100f
C5 z   vss 0.195f
C6 an  vss 0.138f
.ends
