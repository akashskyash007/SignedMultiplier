.subckt noa2a2a2a24_x1 i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa2a2a2a24_x1.ext -        technology: scmos
m00 nq  i7 w1  vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.75555p ps=3.975u
m01 w1  i6 nq  vdd p w=2.19u l=0.13u ad=0.75555p pd=3.975u as=0.58035p ps=2.72u 
m02 w1  i5 w2  vdd p w=2.19u l=0.13u ad=0.75555p pd=3.975u as=0.75555p ps=3.975u
m03 w2  i4 w1  vdd p w=2.19u l=0.13u ad=0.75555p pd=3.975u as=0.75555p ps=3.975u
m04 w3  i3 w2  vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.75555p ps=3.975u
m05 w2  i2 w3  vdd p w=2.19u l=0.13u ad=0.75555p pd=3.975u as=0.58035p ps=2.72u 
m06 w3  i1 vdd vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.93075p ps=5.23u 
m07 vdd i0 w3  vdd p w=2.19u l=0.13u ad=0.93075p pd=5.23u  as=0.58035p ps=2.72u 
m08 w4  i7 vss vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.46325p ps=3.03u 
m09 nq  i6 w4  vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.28885p ps=1.62u 
m10 w5  i5 vss vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.46325p ps=3.03u 
m11 nq  i4 w5  vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.28885p ps=1.62u 
m12 w6  i3 nq  vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.37605p ps=2.325u
m13 vss i2 w6  vss n w=1.09u l=0.13u ad=0.46325p pd=3.03u  as=0.28885p ps=1.62u 
m14 w7  i1 nq  vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.37605p ps=2.325u
m15 vss i0 w7  vss n w=1.09u l=0.13u ad=0.46325p pd=3.03u  as=0.28885p ps=1.62u 
C0  w2 w3  0.073f
C1  nq vdd 0.019f
C2  i5 nq  0.017f
C3  i4 w1  0.005f
C4  i7 i6  0.096f
C5  w2 vdd 0.169f
C6  i4 nq  0.017f
C7  i5 w2  0.005f
C8  i7 vdd 0.010f
C9  nq w4  0.014f
C10 w3 vdd 0.105f
C11 i3 nq  0.017f
C12 i4 w2  0.010f
C13 i1 i0  0.221f
C14 i6 vdd 0.010f
C15 nq w5  0.018f
C16 i2 nq  0.017f
C17 i3 w2  0.014f
C18 i5 vdd 0.010f
C19 nq w6  0.018f
C20 i2 w2  0.005f
C21 i4 vdd 0.010f
C22 i5 i4  0.195f
C23 i2 w3  0.029f
C24 i3 vdd 0.010f
C25 i1 w3  0.041f
C26 w1 nq  0.045f
C27 i2 vdd 0.010f
C28 i4 i3  0.195f
C29 i0 w3  0.012f
C30 w1 w2  0.074f
C31 i1 vdd 0.010f
C32 i7 w1  0.014f
C33 i0 vdd 0.022f
C34 i3 i2  0.195f
C35 i7 nq  0.114f
C36 i6 w1  0.030f
C37 w1 vdd 0.115f
C38 i5 w1  0.023f
C39 i6 nq  0.105f
C40 w7 vss 0.030f
C41 w6 vss 0.026f
C42 w5 vss 0.027f
C43 w4 vss 0.027f
C45 w3 vss 0.061f
C46 w2 vss 0.089f
C47 nq vss 0.488f
C48 w1 vss 0.108f
C49 i0 vss 0.122f
C50 i1 vss 0.135f
C51 i2 vss 0.132f
C52 i3 vss 0.129f
C53 i4 vss 0.118f
C54 i5 vss 0.129f
C55 i6 vss 0.142f
C56 i7 vss 0.157f
.ends
