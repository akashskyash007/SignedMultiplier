* Spice description of vfeed1
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:33
* wsclib 0.13um values
.subckt vfeed1 vdd vss
.ends
