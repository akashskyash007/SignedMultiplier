.subckt nr2v1x3 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2v1x3.ext -        technology: scmos
m00 w1  b z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.37785p  ps=2.58333u
m01 vdd a w1  vdd p w=1.54u l=0.13u ad=0.4081p   pd=2.58333u as=0.19635p  ps=1.795u  
m02 w2  a vdd vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.4081p   ps=2.58333u
m03 z   b w2  vdd p w=1.54u l=0.13u ad=0.37785p  pd=2.58333u as=0.19635p  ps=1.795u  
m04 w3  b z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.37785p  ps=2.58333u
m05 vdd a w3  vdd p w=1.54u l=0.13u ad=0.4081p   pd=2.58333u as=0.19635p  ps=1.795u  
m06 z   b vss vss n w=1.1u  l=0.13u ad=0.231p    pd=1.52u    as=0.488125p ps=2.5375u 
m07 vss a z   vss n w=1.1u  l=0.13u ad=0.488125p pd=2.5375u  as=0.231p    ps=1.52u   
m08 z   b vss vss n w=1.1u  l=0.13u ad=0.231p    pd=1.52u    as=0.488125p ps=2.5375u 
m09 vss a z   vss n w=1.1u  l=0.13u ad=0.488125p pd=2.5375u  as=0.231p    ps=1.52u   
C0  b   z   0.209f
C1  a   z   0.135f
C2  vdd b   0.021f
C3  vdd a   0.032f
C4  a   w2  0.006f
C5  z   w1  0.009f
C6  vdd z   0.071f
C7  a   w3  0.006f
C8  z   w2  0.009f
C9  vdd w1  0.004f
C10 vdd w2  0.004f
C11 vdd w3  0.004f
C12 b   a   0.438f
C13 w3  vss 0.011f
C14 w2  vss 0.009f
C15 w1  vss 0.009f
C16 z   vss 0.470f
C17 a   vss 0.204f
C18 b   vss 0.241f
.ends
