.subckt nd2v0x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v0x2.ext -        technology: scmos
m00 z   b vdd vdd p w=1.32u l=0.13u ad=0.2772p  pd=1.74u  as=0.5313p  ps=3.445u
m01 vdd a z   vdd p w=1.32u l=0.13u ad=0.5313p  pd=3.445u as=0.2772p  ps=1.74u 
m02 w1  b z   vss n w=1.1u  l=0.13u ad=0.14025p pd=1.355u as=0.3278p  ps=2.95u 
m03 vss a w1  vss n w=1.1u  l=0.13u ad=0.5335p  pd=3.17u  as=0.14025p ps=1.355u
C0  b   a   0.134f
C1  b   vdd 0.007f
C2  b   z   0.078f
C3  a   vdd 0.020f
C4  b   w1  0.007f
C5  a   z   0.001f
C6  vdd z   0.086f
C7  w1  vss 0.010f
C8  z   vss 0.217f
C10 a   vss 0.113f
C11 b   vss 0.088f
.ends
