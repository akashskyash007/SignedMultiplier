.subckt vfeed6 vdd vss
*04-JAN-08 SPICE3       file   created      from vfeed6.ext -        technology: scmos
.ends
