* Spice description of bf1v2x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:40:23
* wsclib 0.13um values
.subckt bf1v2x2 a vdd vss z
M01 an    a     vdd   vdd p  L=0.12U  W=0.99U  AS=0.26235P  AD=0.26235P  PS=2.51U   PD=2.51U
M02 an    a     vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M03 vdd   an    z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M04 vss   an    z     vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C3  an    vss   0.471f
C4  a     vss   0.384f
C2  z     vss   0.960f
.ends
