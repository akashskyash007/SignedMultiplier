.subckt iv1v8x1 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v8x1.ext -        technology: scmos
m00 z   a vdd vdd p w=0.825u l=0.13u ad=0.254925p pd=2.4u  as=0.4092p   ps=2.84u
m01 vss a z   vss n w=0.385u l=0.13u ad=0.2563p   pd=2.18u as=0.144375p ps=1.52u
C0 vdd z   0.037f
C1 a   z   0.052f
C2 z   vss 0.140f
C3 a   vss 0.119f
.ends
