* Spice description of aoi21a2bv0x05
* Spice driver version 134999461
* Date  1/01/2008 at 16:36:55
* wsclib 0.13um values
.subckt aoi21a2bv0x05 a1 a2 b vdd vss z
M01 03    a1    vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 vss   a1    sig6  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 vdd   a2n   03    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 sig6  a2n   z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 03    bn    z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M06 z     bn    vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M07 bn    b     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M08 vdd   a2    a2n   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M09 bn    b     vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M10 vss   a2    a2n   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C10 03    vss   0.230f
C8  a1    vss   0.579f
C2  a2n   vss   0.835f
C4  a2    vss   0.619f
C1  bn    vss   0.533f
C5  b     vss   0.631f
C7  z     vss   0.510f
.ends
