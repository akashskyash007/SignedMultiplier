.subckt inv_x2 i nq vdd vss
*05-JAN-08 SPICE3       file   created      from inv_x2.ext -        technology: scmos
m00 nq i vdd vdd p w=1.64u l=0.13u ad=0.697p   pd=4.13u as=1.0666p  ps=5.23u
m01 nq i vss vss n w=1.09u l=0.13u ad=0.46325p pd=3.03u as=0.77235p ps=4.13u
C0 vdd i   0.064f
C1 vdd nq  0.010f
C2 i   nq  0.166f
C3 nq  vss 0.088f
C4 i   vss 0.174f
.ends
