* Sun Dec 16 00:08:09 CET 2007
.subckt xoon21v0x2 a1 a2 b vdd vss z
*SPICE circuit <xoon21v0x2> from XCircuit v3.4 rev 26

m1 an a1 vss vss n w=26u l=2u ad='26u*5u+12p' as='26u*5u+12p' pd='26u*2+14u' ps='26u*2+14u'
m2 an a2 vss vss n w=28u l=2u ad='28u*5u+12p' as='28u*5u+12p' pd='28u*2+14u' ps='28u*2+14u'
m3 n1 a1 vdd vdd p w=70u l=2u ad='70u*5u+12p' as='70u*5u+12p' pd='70u*2+14u' ps='70u*2+14u'
m4 an a2 n1 vdd p w=70u l=2u ad='70u*5u+12p' as='70u*5u+12p' pd='70u*2+14u' ps='70u*2+14u'
m5 z bn an vdd p w=84u l=2u ad='84u*5u+12p' as='84u*5u+12p' pd='84u*2+14u' ps='84u*2+14u'
m6 bn b vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m7 n2 an vss vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m8 z bn n2 vss n w=24u l=2u ad='24u*5u+12p' as='24u*5u+12p' pd='24u*2+14u' ps='24u*2+14u'
m9 bn b vdd vdd p w=47u l=2u ad='47u*5u+12p' as='47u*5u+12p' pd='47u*2+14u' ps='47u*2+14u'
m10 z b an vss n w=18u l=2u ad='18u*5u+12p' as='18u*5u+12p' pd='18u*2+14u' ps='18u*2+14u'
m11 z an bn vdd p w=56u l=2u ad='56u*5u+12p' as='56u*5u+12p' pd='56u*2+14u' ps='56u*2+14u'
.ends
