.subckt mx3_x2 cmd0 cmd1 i0 i1 i2 q vdd vss
*05-JAN-08 SPICE3       file   created      from mx3_x2.ext -        technology: scmos
m00 w1  i2   w2  vdd p w=1.045u l=0.13u ad=0.276925p pd=1.61757u as=0.335426p ps=2.06964u
m01 w3  cmd1 w1  vdd p w=0.99u  l=0.13u ad=0.3663p   pd=2.24836u as=0.26235p  ps=1.53243u
m02 w4  cmd1 vdd vdd p w=0.77u  l=0.13u ad=0.3311p   pd=2.4u     as=0.286694p ps=1.67592u
m03 w5  w4   w3  vdd p w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.38665p  ps=2.37327u
m04 w2  i1   w5  vdd p w=1.045u l=0.13u ad=0.335426p pd=2.06964u as=0.161975p ps=1.355u  
m05 vdd w6   w2  vdd p w=0.99u  l=0.13u ad=0.368607p pd=2.15476u as=0.317772p ps=1.96071u
m06 w7  cmd0 vdd vdd p w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.368607p ps=2.15476u
m07 w3  i0   w7  vdd p w=0.99u  l=0.13u ad=0.3663p   pd=2.24836u as=0.15345p  ps=1.3u    
m08 w4  cmd1 vss vss n w=0.44u  l=0.13u ad=0.1892p   pd=1.74u    as=0.19379p  ps=1.33655u
m09 vdd cmd0 w6  vdd p w=0.77u  l=0.13u ad=0.286694p pd=1.67592u as=0.3311p   ps=2.4u    
m10 q   w3   vdd vdd p w=2.145u l=0.13u ad=0.92235p  pd=5.15u    as=0.798648p ps=4.66864u
m11 w8  i2   w9  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.19u    as=0.24145p  ps=1.70333u
m12 w3  w4   w8  vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u as=0.1749p   ps=1.19u   
m13 w10 cmd1 w3  vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.2959p   ps=2.03333u
m14 w9  i1   w10 vss n w=0.66u  l=0.13u ad=0.24145p  pd=1.70333u as=0.1023p   ps=0.97u   
m15 vss cmd0 w6  vss n w=0.33u  l=0.13u ad=0.145342p pd=1.00241u as=0.1419p   ps=1.52u   
m16 vss cmd0 w9  vss n w=0.66u  l=0.13u ad=0.290685p pd=2.00483u as=0.24145p  ps=1.70333u
m17 w11 w6   vss vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.290685p ps=2.00483u
m18 w3  i0   w11 vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u as=0.1023p   ps=0.97u   
m19 q   w3   vss vss n w=1.1u   l=0.13u ad=0.473p    pd=3.06u    as=0.484474p ps=3.34138u
C0  cmd1 vdd  0.061f
C1  i1   w9   0.007f
C2  vdd  w5   0.010f
C3  i1   cmd0 0.007f
C4  cmd1 w4   0.231f
C5  cmd1 w3   0.023f
C6  w6   w9   0.010f
C7  w2   w1   0.018f
C8  vdd  w7   0.010f
C9  w9   i2   0.007f
C10 w6   cmd0 0.210f
C11 cmd1 w2   0.058f
C12 w2   w5   0.010f
C13 i1   vdd  0.010f
C14 w6   i0   0.165f
C15 w4   i1   0.124f
C16 w9   w8   0.018f
C17 vdd  q    0.034f
C18 i1   w3   0.049f
C19 w6   vdd  0.010f
C20 cmd0 i0   0.219f
C21 vdd  i2   0.010f
C22 w4   i2   0.102f
C23 w9   w10  0.010f
C24 w3   q    0.132f
C25 w6   w3   0.149f
C26 i1   w2   0.007f
C27 cmd0 vdd  0.010f
C28 w4   w9   0.058f
C29 w3   w9   0.057f
C30 i0   vdd  0.010f
C31 cmd0 w3   0.142f
C32 w2   i2   0.007f
C33 cmd1 i1   0.090f
C34 i0   w3   0.043f
C35 w4   vdd  0.010f
C36 cmd1 w6   0.005f
C37 cmd1 i2   0.108f
C38 vdd  w3   0.088f
C39 cmd1 w9   0.007f
C40 w4   w3   0.061f
C41 vdd  w2   0.169f
C42 w4   w2   0.007f
C43 w3   w2   0.085f
C44 vdd  w1   0.017f
C45 i1   w6   0.091f
C46 i1   i2   0.009f
C47 w11  vss  0.012f
C48 w10  vss  0.008f
C49 w8   vss  0.014f
C50 w9   vss  0.218f
C51 q    vss  0.121f
C52 w7   vss  0.007f
C53 w5   vss  0.004f
C54 w1   vss  0.008f
C55 w2   vss  0.059f
C56 w3   vss  0.416f
C58 i0   vss  0.203f
C59 cmd0 vss  0.270f
C60 w6   vss  0.220f
C61 i1   vss  0.136f
C62 w4   vss  0.204f
C63 cmd1 vss  0.308f
C64 i2   vss  0.130f
.ends
