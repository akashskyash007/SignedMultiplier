* Spice description of xnai21v2x05
* Spice driver version 134999461
* Date  1/01/2008 at 17:04:17
* vsclib 0.13um values
.subckt xnai21v2x05 a1 a2 b vdd vss z
M01 a2n   08    z     vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M02 n2    b     vss   vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M03 z     b     vdd   vdd p  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M04 z     a2n   08    vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M05 vss   a2    a2n   vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M06 n1    a2n   n2    vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M07 08    a1    vdd   vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M08 08    a2    z     vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M09 vdd   a2    a2n   vdd p  L=0.12U  W=1.155U AS=0.306075P AD=0.306075P PS=2.84U   PD=2.84U
M10 z     08    n1    vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
M11 n2    a1    08    vss n  L=0.12U  W=0.715U AS=0.189475P AD=0.189475P PS=1.96U   PD=1.96U
C7  08    vss   0.769f
C9  a1    vss   0.754f
C2  a2n   vss   0.929f
C4  a2    vss   0.953f
C5  b     vss   0.364f
C1  n2    vss   0.231f
C6  z     vss   0.673f
.ends
