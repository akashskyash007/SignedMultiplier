.subckt oai22v0x05 a1 a2 b1 b2 vdd vss z
*01-JAN-08 SPICE3       file   created      from oai22v0x05.ext -        technology: scmos
m00 w1  b1 vdd vdd p w=0.88u  l=0.13u ad=0.1364p   pd=1.19u   as=0.431338p ps=2.895u 
m01 z   b2 w1  vdd p w=0.88u  l=0.13u ad=0.1848p   pd=1.3u    as=0.1364p   ps=1.19u  
m02 w2  a2 z   vdd p w=0.88u  l=0.13u ad=0.1364p   pd=1.19u   as=0.1848p   ps=1.3u   
m03 vdd a1 w2  vdd p w=0.88u  l=0.13u ad=0.431338p pd=2.895u  as=0.1364p   ps=1.19u  
m04 n3  b2 z   vss n w=0.385u l=0.13u ad=0.112613p pd=1.1625u as=0.133788p ps=1.245u 
m05 vss a2 n3  vss n w=0.385u l=0.13u ad=0.221513p pd=1.795u  as=0.112613p ps=1.1625u
m06 z   b1 n3  vss n w=0.385u l=0.13u ad=0.133788p pd=1.245u  as=0.112613p ps=1.1625u
m07 n3  a1 vss vss n w=0.385u l=0.13u ad=0.112613p pd=1.1625u as=0.221513p ps=1.795u 
C0  a1  z   0.016f
C1  b2  n3  0.005f
C2  vdd b1  0.006f
C3  a2  n3  0.063f
C4  a1  w2  0.022f
C5  w1  z   0.010f
C6  vdd b2  0.006f
C7  a1  n3  0.006f
C8  vdd a2  0.006f
C9  vdd a1  0.034f
C10 b1  b2  0.116f
C11 z   n3  0.082f
C12 b1  a2  0.009f
C13 vdd w1  0.003f
C14 vdd z   0.115f
C15 b2  a2  0.082f
C16 vdd w2  0.003f
C17 b2  a1  0.006f
C18 b1  z   0.109f
C19 b2  w1  0.005f
C20 a2  a1  0.090f
C21 b2  z   0.022f
C22 b1  n3  0.006f
C23 n3  vss 0.244f
C24 w2  vss 0.007f
C25 z   vss 0.172f
C26 w1  vss 0.006f
C27 a1  vss 0.116f
C28 a2  vss 0.117f
C29 b2  vss 0.094f
C30 b1  vss 0.107f
.ends
