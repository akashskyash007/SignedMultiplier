.subckt cgi2v0x05 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from cgi2v0x05.ext -        technology: scmos
m00 vdd a n1  vdd p w=0.88u  l=0.13u ad=0.358233p  pd=2.84u    as=0.22715p   ps=1.70333u
m01 w1  a vdd vdd p w=0.88u  l=0.13u ad=0.1122p    pd=1.135u   as=0.358233p  ps=2.84u   
m02 z   b w1  vdd p w=0.88u  l=0.13u ad=0.1848p    pd=1.3u     as=0.1122p    ps=1.135u  
m03 n1  c z   vdd p w=0.88u  l=0.13u ad=0.22715p   pd=1.70333u as=0.1848p    ps=1.3u    
m04 vdd b n1  vdd p w=0.88u  l=0.13u ad=0.358233p  pd=2.84u    as=0.22715p   ps=1.70333u
m05 w2  a vss vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u    as=0.23815p   ps=2.18u   
m06 z   b w2  vss n w=0.385u l=0.13u ad=0.08085p   pd=0.805u   as=0.0490875p ps=0.64u   
m07 n3  c z   vss n w=0.385u l=0.13u ad=0.102025p  pd=1.04333u as=0.08085p   ps=0.805u  
m08 vss b n3  vss n w=0.385u l=0.13u ad=0.23815p   pd=2.18u    as=0.102025p  ps=1.04333u
m09 vss a n3  vss n w=0.385u l=0.13u ad=0.23815p   pd=2.18u    as=0.102025p  ps=1.04333u
C0  z   w2  0.007f
C1  vdd n1  0.126f
C2  b   a   0.094f
C3  z   n3  0.073f
C4  b   c   0.167f
C5  vdd z   0.022f
C6  b   n1  0.033f
C7  a   c   0.006f
C8  a   n1  0.021f
C9  b   z   0.014f
C10 c   n1  0.007f
C11 a   z   0.063f
C12 b   n3  0.005f
C13 c   z   0.106f
C14 n1  z   0.133f
C15 a   n3  0.053f
C16 vdd b   0.047f
C17 c   n3  0.005f
C18 w1  z   0.014f
C19 n3  vss 0.225f
C20 z   vss 0.090f
C21 w1  vss 0.004f
C22 n1  vss 0.100f
C23 c   vss 0.083f
C24 a   vss 0.177f
C25 b   vss 0.177f
.ends
