.subckt cgi2_x05 a b c vdd vss z
*04-JAN-08 SPICE3       file   created      from cgi2_x05.ext -        technology: scmos
m00 vdd a n2  vdd p w=1.1u   l=0.13u ad=0.352p    pd=2.10667u as=0.33385p  ps=2.10667u
m01 w1  a vdd vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u    as=0.352p    ps=2.10667u
m02 z   b w1  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.1705p   ps=1.41u   
m03 n2  c z   vdd p w=1.1u   l=0.13u ad=0.33385p  pd=2.10667u as=0.2915p   ps=1.63u   
m04 vdd b n2  vdd p w=1.1u   l=0.13u ad=0.352p    pd=2.10667u as=0.33385p  ps=2.10667u
m05 vss a n4  vss n w=0.495u l=0.13u ad=0.2673p   pd=1.96u    as=0.149325p ps=1.3u    
m06 w2  a vss vss n w=0.495u l=0.13u ad=0.076725p pd=0.805u   as=0.2673p   ps=1.96u   
m07 z   b w2  vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u   as=0.076725p ps=0.805u  
m08 n4  c z   vss n w=0.495u l=0.13u ad=0.149325p pd=1.3u     as=0.131175p ps=1.025u  
m09 vss b n4  vss n w=0.495u l=0.13u ad=0.2673p   pd=1.96u    as=0.149325p ps=1.3u    
C0  w3  c   0.001f
C1  w4  b   0.015f
C2  c   n4  0.004f
C3  n2  z   0.056f
C4  vdd a   0.004f
C5  w3  n2  0.043f
C6  w4  c   0.018f
C7  w1  z   0.002f
C8  vdd b   0.006f
C9  w5  w4  0.166f
C10 w3  w1  0.002f
C11 w4  n2  0.022f
C12 vdd c   0.016f
C13 w3  z   0.005f
C14 w4  w1  0.005f
C15 w6  z   0.009f
C16 z   n4  0.058f
C17 vdd n2  0.146f
C18 a   b   0.117f
C19 w4  z   0.023f
C20 z   w2  0.014f
C21 w3  w4  0.166f
C22 w5  a   0.013f
C23 w6  w4  0.166f
C24 w4  n4  0.060f
C25 a   n2  0.028f
C26 b   c   0.243f
C27 w5  b   0.010f
C28 w3  vdd 0.025f
C29 w4  w2  0.002f
C30 b   n2  0.007f
C31 w5  c   0.011f
C32 w4  vdd 0.044f
C33 a   z   0.019f
C34 c   n2  0.056f
C35 w3  a   0.005f
C36 w6  a   0.013f
C37 a   n4  0.010f
C38 b   z   0.061f
C39 w3  b   0.004f
C40 w4  a   0.019f
C41 w6  b   0.059f
C42 c   z   0.041f
C43 b   n4  0.019f
C44 n2  w1  0.029f
C45 w5  z   0.030f
C46 w4  vss 1.000f
C47 w6  vss 0.171f
C48 w5  vss 0.175f
C49 w3  vss 0.159f
C50 n4  vss 0.203f
C51 z   vss 0.037f
C52 n2  vss 0.002f
C53 c   vss 0.081f
C54 b   vss 0.167f
C55 a   vss 0.172f
.ends
