.subckt bf1v2x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v2x2.ext -        technology: scmos
m00 vdd an z   vdd p w=1.54u  l=0.13u ad=0.463339p pd=2.52u    as=0.48675p  ps=3.83u   
m01 an  a  vdd vdd p w=0.99u  l=0.13u ad=0.29865p  pd=2.73u    as=0.297861p ps=1.62u   
m02 vss an z   vss n w=0.77u  l=0.13u ad=0.23167p  pd=1.58261u as=0.28875p  ps=2.29u   
m03 an  a  vss vss n w=0.495u l=0.13u ad=0.167475p pd=1.74u    as=0.14893p  ps=1.01739u
C0 vdd an  0.039f
C1 vdd z   0.054f
C2 an  z   0.135f
C3 an  a   0.155f
C4 a   vss 0.101f
C5 z   vss 0.193f
C6 an  vss 0.140f
.ends
