.subckt oai21bv0x05 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from oai21bv0x05.ext -        technology: scmos
m00 z   bn vdd vdd p w=0.44u  l=0.13u ad=0.100467p pd=0.866667u as=0.175676p ps=1.25412u
m01 w1  a2 z   vdd p w=0.88u  l=0.13u ad=0.1122p   pd=1.135u    as=0.200933p ps=1.73333u
m02 vdd a1 w1  vdd p w=0.88u  l=0.13u ad=0.351353p pd=2.50824u  as=0.1122p   ps=1.135u  
m03 bn  b  vdd vdd p w=0.55u  l=0.13u ad=0.18205p  pd=1.85u     as=0.219596p ps=1.56765u
m04 n1  bn z   vss n w=0.385u l=0.13u ad=0.102025p pd=1.04333u  as=0.144375p ps=1.52u   
m05 vss a2 n1  vss n w=0.385u l=0.13u ad=0.21637p  pd=1.75u     as=0.102025p ps=1.04333u
m06 vss b  bn  vss n w=0.33u  l=0.13u ad=0.18546p  pd=1.5u      as=0.12375p  ps=1.41u   
m07 n1  a1 vss vss n w=0.385u l=0.13u ad=0.102025p pd=1.04333u  as=0.21637p  ps=1.75u   
C0  bn  a1  0.124f
C1  bn  z   0.082f
C2  a2  a1  0.169f
C3  bn  w1  0.008f
C4  a2  z   0.007f
C5  a1  z   0.050f
C6  bn  b   0.041f
C7  a2  n1  0.019f
C8  a1  b   0.021f
C9  a1  n1  0.009f
C10 vdd bn  0.038f
C11 z   n1  0.026f
C12 vdd a2  0.005f
C13 vdd a1  0.005f
C14 vdd z   0.087f
C15 bn  a2  0.106f
C16 n1  vss 0.144f
C17 b   vss 0.121f
C18 w1  vss 0.005f
C19 z   vss 0.199f
C20 a1  vss 0.118f
C21 a2  vss 0.110f
C22 bn  vss 0.163f
.ends
