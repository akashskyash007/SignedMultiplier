* Spice description of vfeed8
* Spice driver version 134999461
* Date  1/01/2008 at 17:03:09
* vsclib 0.13um values
.subckt vfeed8 vdd vss
.ends
