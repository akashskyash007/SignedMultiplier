.subckt rowend_x0 vdd vss
*04-JAN-08 SPICE3       file   created      from rowend_x0.ext -        technology: scmos
C0 vdd w1  0.005f
C1 w2  w1  0.166f
C2 w3  w1  0.166f
C3 w4  w1  0.166f
C4 w1  vss 1.089f
C5 w4  vss 0.196f
C6 w3  vss 0.196f
C7 w2  vss 0.196f
.ends
