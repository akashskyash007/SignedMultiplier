.subckt cgi2a_x1 a b c vdd vss z
*04-JAN-08 SPICE3       file   created      from cgi2a_x1.ext -        technology: scmos
m00 vdd b  n2  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.610775p ps=3.5u  
m01 w1  b  vdd vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=0.568425p ps=2.675u
m02 z   an w1  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.332475p ps=2.455u
m03 n2  c  z   vdd p w=2.145u l=0.13u ad=0.610775p pd=3.5u   as=0.568425p ps=2.675u
m04 vdd an n2  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.610775p ps=3.5u  
m05 an  a  vdd vdd p w=2.145u l=0.13u ad=0.622875p pd=5.15u  as=0.568425p ps=2.675u
m06 vss b  n4  vss n w=0.99u  l=0.13u ad=0.289575p pd=1.685u as=0.3047p   ps=1.96u 
m07 w2  b  vss vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u   as=0.289575p ps=1.685u
m08 z   an w2  vss n w=0.99u  l=0.13u ad=0.26235p  pd=1.52u  as=0.15345p  ps=1.3u  
m09 n4  c  z   vss n w=0.99u  l=0.13u ad=0.3047p   pd=1.96u  as=0.26235p  ps=1.52u 
m10 vss an n4  vss n w=0.99u  l=0.13u ad=0.289575p pd=1.685u as=0.3047p   ps=1.96u 
m11 an  a  vss vss n w=0.99u  l=0.13u ad=0.3894p   pd=2.84u  as=0.289575p ps=1.685u
C0  n4  w2  0.020f
C1  c   vdd 0.010f
C2  b   n4  0.029f
C3  an  z   0.015f
C4  a   vdd 0.069f
C5  an  n4  0.023f
C6  c   z   0.096f
C7  n2  vdd 0.172f
C8  c   n4  0.007f
C9  n2  w1  0.029f
C10 n2  z   0.024f
C11 vdd w1  0.010f
C12 b   an  0.151f
C13 vdd z   0.017f
C14 w1  z   0.009f
C15 an  c   0.202f
C16 b   n2  0.036f
C17 an  a   0.152f
C18 z   n4  0.075f
C19 an  n2  0.007f
C20 b   vdd 0.020f
C21 c   a   0.076f
C22 c   n2  0.103f
C23 an  vdd 0.029f
C24 w2  vss 0.005f
C25 n4  vss 0.237f
C26 z   vss 0.089f
C27 w1  vss 0.009f
C29 n2  vss 0.098f
C30 a   vss 0.101f
C31 c   vss 0.111f
C32 an  vss 0.346f
C33 b   vss 0.191f
.ends
