.subckt bf1_w2 a vdd vss z
*04-JAN-08 SPICE3       file   created      from bf1_w2.ext -        technology: scmos
m00 vdd an z   vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u  as=0.6809p   ps=5.04u 
m01 an  a  vdd vdd p w=2.09u  l=0.13u ad=0.6809p   pd=5.04u  as=0.55385p  ps=2.62u 
m02 vss an z   vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u as=0.403975p ps=2.95u 
m03 an  a  vss vss n w=1.045u l=0.13u ad=0.403975p pd=2.95u  as=0.276925p ps=1.575u
C0 z  vdd 0.008f
C1 an a   0.215f
C2 an z   0.111f
C3 an vdd 0.083f
C4 a  vdd 0.010f
C6 z  vss 0.111f
C7 a  vss 0.105f
C8 an vss 0.218f
.ends
