* Spice description of bf1_y1
* Spice driver version 134999461
* Date  4/01/2008 at 18:54:47
* vsxlib 0.13um values
.subckt bf1_y1 a vdd vss z
M1a 2z    a     vdd   vdd p  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M1z vdd   2z    z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2a vss   a     2z    vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M2z z     2z    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C4  2z    vss   0.869f
C3  a     vss   0.714f
C2  z     vss   0.506f
.ends
