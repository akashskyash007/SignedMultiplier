.subckt nxr2_x1 i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nxr2_x1.ext -        technology: scmos
m00 vdd i0 w1  vdd p w=1.09u l=0.13u ad=0.347338p pd=1.80781u as=0.46325p  ps=3.03u   
m01 w2  i0 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.697862p ps=3.6322u 
m02 nq  i1 w2  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.58035p  ps=2.72u   
m03 w2  w1 nq  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.58035p  ps=2.72u   
m04 vdd w3 w2  vdd p w=2.19u l=0.13u ad=0.697862p pd=3.6322u  as=0.58035p  ps=2.72u   
m05 w3  i1 vdd vdd p w=1.09u l=0.13u ad=0.58315p  pd=3.25u    as=0.347338p ps=1.80781u
m06 vss i0 w1  vss n w=0.54u l=0.13u ad=0.172253p pd=1.07337u as=0.2295p   ps=1.93u   
m07 w4  i0 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.347697p ps=2.16663u
m08 nq  w3 w4  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.28885p  ps=1.62u   
m09 w5  w1 nq  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.28885p  ps=1.62u   
m10 vss i1 w5  vss n w=1.09u l=0.13u ad=0.347697p pd=2.16663u as=0.28885p  ps=1.62u   
m11 w3  i1 vss vss n w=0.54u l=0.13u ad=0.2889p   pd=2.15u    as=0.172253p ps=1.07337u
C0  nq  w4  0.018f
C1  vdd w3  0.021f
C2  i0  i1  0.047f
C3  vdd w2  0.103f
C4  i0  w1  0.138f
C5  vdd nq  0.019f
C6  i0  w3  0.027f
C7  i1  w1  0.108f
C8  i0  w2  0.010f
C9  i1  w3  0.261f
C10 i0  nq  0.140f
C11 i1  w2  0.014f
C12 w1  w3  0.132f
C13 i1  nq  0.017f
C14 w1  w2  0.005f
C15 w1  nq  0.007f
C16 w3  nq  0.032f
C17 vdd i0  0.075f
C18 w2  nq  0.095f
C19 vdd i1  0.050f
C20 vdd w1  0.021f
C21 w5  vss 0.030f
C22 w4  vss 0.027f
C23 nq  vss 0.169f
C24 w2  vss 0.065f
C25 w3  vss 0.247f
C26 w1  vss 0.332f
C27 i1  vss 0.259f
C28 i0  vss 0.229f
.ends
