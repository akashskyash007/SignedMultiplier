.subckt nd2abv0x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2abv0x2.ext -        technology: scmos
m00 vdd b  bn  vdd p w=0.99u  l=0.13u ad=0.302539p pd=1.70357u as=0.341p    ps=2.73u   
m01 z   bn vdd vdd p w=1.32u  l=0.13u ad=0.2772p   pd=1.74u    as=0.403386p ps=2.27143u
m02 vdd an z   vdd p w=1.32u  l=0.13u ad=0.403386p pd=2.27143u as=0.2772p   ps=1.74u   
m03 an  a  vdd vdd p w=0.99u  l=0.13u ad=0.29865p  pd=2.73u    as=0.302539p ps=1.70357u
m04 vss b  bn  vss n w=0.495u l=0.13u ad=0.16843p  pd=1.31447u as=0.167475p ps=1.74u   
m05 w1  bn z   vss n w=1.1u   l=0.13u ad=0.14025p  pd=1.355u   as=0.3278p   ps=2.95u   
m06 vss an w1  vss n w=1.1u   l=0.13u ad=0.37429p  pd=2.92105u as=0.14025p  ps=1.355u  
m07 an  a  vss vss n w=0.495u l=0.13u ad=0.167475p pd=1.74u    as=0.16843p  ps=1.31447u
C0  bn  an  0.107f
C1  vdd z   0.031f
C2  bn  b   0.105f
C3  an  a   0.162f
C4  bn  z   0.053f
C5  an  z   0.010f
C6  a   z   0.023f
C7  b   z   0.069f
C8  b   w1  0.004f
C9  vdd bn  0.006f
C10 vdd an  0.016f
C11 vdd a   0.051f
C12 w1  vss 0.011f
C13 z   vss 0.063f
C14 b   vss 0.166f
C15 a   vss 0.101f
C16 an  vss 0.160f
C17 bn  vss 0.253f
.ends
