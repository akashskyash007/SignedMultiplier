* Spice description of nr2a_x05
* Spice driver version 134999461
* Date  4/01/2008 at 19:06:46
* vxlib 0.13um values
.subckt nr2a_x05 a b vdd vss z
M1a an    a     vdd   vdd p  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M1z vdd   an    sig4  vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M2a vss   a     an    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M2z sig4  b     z     vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M3z z     an    vss   vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
M4z vss   b     z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C3  an    vss   0.873f
C6  a     vss   0.847f
C7  b     vss   0.927f
C1  z     vss   0.701f
.ends
