* Spice description of nr2a_x1
* Spice driver version 134999461
* Date  4/01/2008 at 19:07:02
* vxlib 0.13um values
.subckt nr2a_x1 a b vdd vss z
M1a sig2  a     vdd   vdd p  L=0.12U  W=1.21U  AS=0.32065P  AD=0.32065P  PS=2.95U   PD=2.95U
M1z vdd   sig2  sig4  vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2a vss   a     sig2  vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
M2z sig4  b     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M3z z     sig2  vss   vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
M4z vss   b     z     vss n  L=0.12U  W=0.605U AS=0.160325P AD=0.160325P PS=1.74U   PD=1.74U
C6  a     vss   0.831f
C7  b     vss   0.886f
C2  sig2  vss   0.818f
C3  z     vss   0.701f
.ends
