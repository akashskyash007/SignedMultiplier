.subckt nr2a_x05 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2a_x05.ext -        technology: scmos
m00 w1  b  z   vdd p w=1.21u  l=0.13u ad=0.18755p  pd=1.52u    as=0.4477p   ps=3.28u   
m01 vdd an w1  vdd p w=1.21u  l=0.13u ad=0.421328p pd=2.08718u as=0.18755p  ps=1.52u   
m02 an  a  vdd vdd p w=0.935u l=0.13u ad=0.374825p pd=2.73u    as=0.325572p ps=1.61282u
m03 z   b  vss vss n w=0.33u  l=0.13u ad=0.08745p  pd=0.86u    as=0.173879p ps=1.36571u
m04 vss an z   vss n w=0.33u  l=0.13u ad=0.173879p pd=1.36571u as=0.08745p  ps=0.86u   
m05 an  a  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.260818p ps=2.04857u
C0  vdd an  0.005f
C1  b   an  0.160f
C2  b   z   0.099f
C3  vdd a   0.049f
C4  b   a   0.031f
C5  an  a   0.145f
C6  z   a   0.041f
C7  w1  a   0.033f
C8  a   vss 0.134f
C9  w1  vss 0.004f
C10 z   vss 0.180f
C11 an  vss 0.200f
C12 b   vss 0.158f
.ends
