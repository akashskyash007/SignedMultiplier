.subckt halfadder_x4 a b cout sout vdd vss
*05-JAN-08 SPICE3       file   created      from halfadder_x4.ext -        technology: scmos
m00 cout w1 vdd  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.864224p ps=4.98175u
m01 vdd  w1 cout vdd p w=2.145u l=0.13u ad=0.864224p pd=4.98175u as=0.568425p ps=2.675u  
m02 w1   a  vdd  vdd p w=0.99u  l=0.13u ad=0.266888p pd=1.575u   as=0.398872p ps=2.29927u
m03 vdd  b  w1   vdd p w=0.99u  l=0.13u ad=0.398872p pd=2.29927u as=0.266888p ps=1.575u  
m04 vdd  b  w2   vdd p w=0.88u  l=0.13u ad=0.354553p pd=2.0438u  as=0.3784p   ps=2.62u   
m05 w3   b  vdd  vdd p w=1.21u  l=0.13u ad=0.32065p  pd=1.74u    as=0.487511p ps=2.81022u
m06 w4   a  w3   vdd p w=1.21u  l=0.13u ad=0.325188p pd=1.795u   as=0.32065p  ps=1.74u   
m07 w3   w2 w4   vdd p w=1.21u  l=0.13u ad=0.32065p  pd=1.74u    as=0.325188p ps=1.795u  
m08 vdd  w5 w3   vdd p w=1.21u  l=0.13u ad=0.487511p pd=2.81022u as=0.32065p  ps=1.74u   
m09 w5   a  vdd  vdd p w=1.21u  l=0.13u ad=0.5687p   pd=3.61u    as=0.487511p ps=2.81022u
m10 sout w4 vdd  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.864224p ps=4.98175u
m11 vdd  w4 sout vdd p w=2.145u l=0.13u ad=0.864224p pd=4.98175u as=0.568425p ps=2.675u  
m12 cout w1 vss  vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.416024p ps=2.8516u 
m13 vss  w1 cout vss n w=1.045u l=0.13u ad=0.416024p pd=2.8516u  as=0.276925p ps=1.575u  
m14 w6   a  vss  vss n w=0.495u l=0.13u ad=0.14893p  pd=1.01739u as=0.197064p ps=1.35076u
m15 w1   b  w6   vss n w=0.77u  l=0.13u ad=0.3311p   pd=2.4u     as=0.23167p  ps=1.58261u
m16 vss  b  w2   vss n w=0.44u  l=0.13u ad=0.175168p pd=1.20067u as=0.180125p ps=1.74u   
m17 w7   b  vss  vss n w=0.495u l=0.13u ad=0.139343p pd=1.0215u  as=0.197064p ps=1.35076u
m18 w4   w5 w7   vss n w=0.605u l=0.13u ad=0.160325p pd=1.13826u as=0.170308p ps=1.2485u 
m19 w8   w2 w4   vss n w=0.66u  l=0.13u ad=0.190457p pd=1.36u    as=0.1749p   ps=1.24174u
m20 vss  a  w8   vss n w=0.495u l=0.13u ad=0.197064p pd=1.35076u as=0.142843p ps=1.02u   
m21 w5   a  vss  vss n w=0.44u  l=0.13u ad=0.38885p  pd=2.95u    as=0.175168p ps=1.20067u
m22 sout w4 vss  vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.416024p ps=2.8516u 
m23 vss  w4 sout vss n w=1.045u l=0.13u ad=0.416024p pd=2.8516u  as=0.276925p ps=1.575u  
C0  w3   w4   0.087f
C1  w2   w5   0.116f
C2  w1   cout 0.020f
C3  vdd  b    0.058f
C4  w7   w4   0.020f
C5  w1   a    0.271f
C6  w8   w4   0.018f
C7  w4   w5   0.137f
C8  sout w4   0.085f
C9  cout a    0.171f
C10 w1   b    0.128f
C11 w6   w1   0.025f
C12 w1   w2   0.009f
C13 vdd  w4   0.020f
C14 a    b    0.176f
C15 sout vdd  0.127f
C16 a    w2   0.083f
C17 a    w3   0.101f
C18 b    w2   0.154f
C19 b    w3   0.012f
C20 a    w4   0.069f
C21 vdd  w1   0.020f
C22 b    w4   0.114f
C23 w2   w3   0.007f
C24 a    w5   0.232f
C25 vdd  cout 0.086f
C26 w2   w4   0.014f
C27 b    w5   0.018f
C28 vdd  a    0.390f
C29 w8   vss  0.007f
C30 w7   vss  0.007f
C31 w6   vss  0.005f
C32 sout vss  0.145f
C33 w5   vss  0.224f
C34 w4   vss  0.589f
C35 w3   vss  0.045f
C36 w2   vss  0.234f
C37 b    vss  0.364f
C38 a    vss  0.554f
C39 cout vss  0.145f
C40 w1   vss  0.370f
.ends
