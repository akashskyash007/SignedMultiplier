.subckt vsstie vdd vss z
*01-JAN-08 SPICE3       file   created      from vsstie.ext -        technology: scmos
m00 z   vdd vdd vdd p w=0.99u l=0.13u ad=0.4257p pd=2.84u as=0.73425p ps=4.27u
m01 vss vdd z   vss n w=1.1u  l=0.13u ad=0.473p  pd=3.06u as=0.5335p  ps=3.17u
C0 vdd z   0.103f
C1 z   vss 0.209f
.ends
