.subckt nmx3_x1 cmd0 cmd1 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nmx3_x1.ext -        technology: scmos
m00 w1  i2   w2  vdd p w=1.045u l=0.13u ad=0.276925p pd=1.61757u as=0.3344p   ps=2.03333u
m01 nq  cmd1 w1  vdd p w=0.99u  l=0.13u ad=0.367361p pd=2.24357u as=0.26235p  ps=1.53243u
m02 w3  cmd1 vdd vdd p w=0.77u  l=0.13u ad=0.3311p   pd=2.4u     as=0.3619p   ps=2.31636u
m03 w4  w3   nq  vdd p w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.38777p  ps=2.36821u
m04 w2  i1   w4  vdd p w=1.045u l=0.13u ad=0.3344p   pd=2.03333u as=0.161975p ps=1.355u  
m05 vdd w5   w2  vdd p w=1.045u l=0.13u ad=0.49115p  pd=3.14364u as=0.3344p   ps=2.03333u
m06 w6  cmd0 vdd vdd p w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.49115p  ps=3.14364u
m07 nq  i0   w6  vdd p w=1.045u l=0.13u ad=0.38777p  pd=2.36821u as=0.161975p ps=1.355u  
m08 w3  cmd1 vss vss n w=0.44u  l=0.13u ad=0.1892p   pd=1.74u    as=0.27027p  ps=1.942u  
m09 vdd cmd0 w5  vdd p w=0.77u  l=0.13u ad=0.3619p   pd=2.31636u as=0.3311p   ps=2.4u    
m10 w7  i2   w8  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.19u    as=0.24145p  ps=1.70333u
m11 nq  w3   w7  vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u as=0.1749p   ps=1.19u   
m12 w9  cmd1 nq  vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.2959p   ps=2.03333u
m13 w8  i1   w9  vss n w=0.66u  l=0.13u ad=0.24145p  pd=1.70333u as=0.1023p   ps=0.97u   
m14 vss cmd0 w5  vss n w=0.44u  l=0.13u ad=0.27027p  pd=1.942u   as=0.1892p   ps=1.74u   
m15 vss cmd0 w8  vss n w=0.66u  l=0.13u ad=0.405405p pd=2.913u   as=0.24145p  ps=1.70333u
m16 w10 w5   vss vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.405405p ps=2.913u  
m17 nq  i0   w10 vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u as=0.1023p   ps=0.97u   
C0  i1   w2   0.007f
C1  w3   i1   0.124f
C2  i0   vdd  0.010f
C3  w2   cmd1 0.058f
C4  w3   cmd1 0.232f
C5  nq   w8   0.030f
C6  w5   nq   0.141f
C7  i1   nq   0.073f
C8  cmd0 nq   0.098f
C9  vdd  w2   0.169f
C10 w3   vdd  0.010f
C11 nq   cmd1 0.028f
C12 i0   nq   0.043f
C13 vdd  w1   0.017f
C14 w3   w2   0.007f
C15 w2   w1   0.018f
C16 vdd  nq   0.107f
C17 w5   w8   0.010f
C18 w2   nq   0.085f
C19 vdd  w4   0.010f
C20 w3   nq   0.058f
C21 w8   i2   0.007f
C22 w8   w7   0.018f
C23 i1   w8   0.007f
C24 w2   w4   0.010f
C25 vdd  w6   0.010f
C26 i1   w5   0.092f
C27 w8   cmd1 0.007f
C28 w5   cmd0 0.209f
C29 i1   i2   0.009f
C30 w5   cmd1 0.005f
C31 i2   cmd1 0.108f
C32 w8   w9   0.010f
C33 i1   cmd0 0.007f
C34 w5   i0   0.165f
C35 i1   cmd1 0.090f
C36 w5   vdd  0.010f
C37 cmd0 i0   0.218f
C38 vdd  i2   0.010f
C39 i1   vdd  0.010f
C40 w3   w8   0.058f
C41 cmd0 vdd  0.010f
C42 w2   i2   0.007f
C43 vdd  cmd1 0.061f
C44 w3   i2   0.102f
C45 w10  vss  0.012f
C46 w9   vss  0.008f
C47 w7   vss  0.014f
C48 w8   vss  0.218f
C49 w6   vss  0.007f
C50 w4   vss  0.004f
C51 nq   vss  0.355f
C52 w1   vss  0.008f
C53 w2   vss  0.059f
C55 i0   vss  0.201f
C56 cmd0 vss  0.265f
C57 w5   vss  0.216f
C58 i1   vss  0.136f
C59 w3   vss  0.205f
C60 cmd1 vss  0.306f
C61 i2   vss  0.130f
.ends
