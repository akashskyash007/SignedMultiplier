.subckt an2_x2 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from an2_x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=2.09u  l=0.13u ad=0.702763p pd=3.82159u as=0.6809p   ps=5.04u   
m01 zn  a  vdd vdd p w=1.375u l=0.13u ad=0.364375p pd=1.905u   as=0.462344p ps=2.5142u 
m02 vdd b  zn  vdd p w=1.375u l=0.13u ad=0.462344p pd=2.5142u  as=0.364375p ps=1.905u  
m03 vss zn z   vss n w=1.045u l=0.13u ad=0.345895p pd=1.70525u as=0.403975p ps=2.95u   
m04 w1  a  vss vss n w=1.155u l=0.13u ad=0.179025p pd=1.465u   as=0.382305p ps=1.88475u
m05 zn  b  w1  vss n w=1.155u l=0.13u ad=0.433125p pd=3.17u    as=0.179025p ps=1.465u  
C0  zn  a   0.187f
C1  zn  b   0.077f
C2  zn  w1  0.010f
C3  z   b   0.016f
C4  a   b   0.155f
C5  a   w1  0.004f
C6  vdd zn  0.031f
C7  vdd z   0.036f
C8  vdd a   0.002f
C9  zn  z   0.119f
C10 vdd b   0.020f
C11 w1  vss 0.007f
C12 b   vss 0.092f
C13 a   vss 0.116f
C14 z   vss 0.081f
C15 zn  vss 0.227f
.ends
