.subckt nao22_x1 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nao22_x1.ext -        technology: scmos
m00 w1  i0 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u as=0.93075p  ps=5.23u
m01 nq  i1 w1  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u as=0.58035p  ps=2.72u
m02 vdd i2 nq  vdd p w=2.19u l=0.13u ad=0.93075p  pd=5.23u as=0.58035p  ps=2.72u
m03 nq  i0 w2  vss n w=1.09u l=0.13u ad=0.35925p  pd=2.06u as=0.346983p ps=2.09u
m04 w2  i1 nq  vss n w=1.09u l=0.13u ad=0.346983p pd=2.09u as=0.35925p  ps=2.06u
m05 vss i2 w2  vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u as=0.346983p ps=2.09u
C0  vdd w1  0.019f
C1  i0  i1  0.221f
C2  vdd nq  0.029f
C3  i1  i2  0.096f
C4  i1  w1  0.052f
C5  i1  nq  0.132f
C6  i0  w2  0.005f
C7  i1  w2  0.005f
C8  i2  nq  0.140f
C9  i2  w2  0.010f
C10 vdd i0  0.052f
C11 nq  w2  0.051f
C12 vdd i1  0.021f
C13 vdd i2  0.113f
C14 w2  vss 0.139f
C15 nq  vss 0.122f
C16 w1  vss 0.015f
C17 i2  vss 0.210f
C18 i1  vss 0.133f
C19 i0  vss 0.132f
.ends
