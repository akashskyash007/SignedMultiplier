.subckt mxi2v2x1 a0 a1 s vdd vss z
*10-JAN-08 SPICE3       file   created      from mxi2v2x1.ext -        technology: scmos
m00 vdd a1  w1  vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 w2  a0  vdd vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 z   w3  w1  vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m03 w2  s   z   vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m04 vdd s   w3  vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m05 w4  vdd vdd vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m06 vss a1  w1  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m07 w2  a0  vss vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
m08 z   w3  w2  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m09 w1  s   z   vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
m10 vss s   w3  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m11 w5  vdd vss vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0  vdd z   0.010f
C1  a1  a0  0.089f
C2  w1  a0  0.129f
C3  vdd s   0.103f
C4  w1  w3  0.034f
C5  w1  z   0.031f
C6  a0  w3  0.050f
C7  w1  s   0.030f
C8  w3  z   0.095f
C9  w1  w2  0.140f
C10 a0  w2  0.110f
C11 w3  s   0.225f
C12 vdd a1  0.007f
C13 z   s   0.091f
C14 w3  w2  0.208f
C15 vdd w1  0.070f
C16 z   w2  0.049f
C17 vdd a0  0.007f
C18 s   w2  0.011f
C19 vdd w3  0.062f
C20 a1  w1  0.132f
C21 w5  vss 0.014f
C22 w4  vss 0.019f
C23 w2  vss 0.132f
C24 s   vss 0.295f
C25 z   vss 0.072f
C26 w3  vss 0.271f
C27 a0  vss 0.149f
C28 w1  vss 0.434f
C29 a1  vss 0.153f
.ends
