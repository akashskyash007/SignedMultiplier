.subckt bf1v0x12 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v0x12.ext -        technology: scmos
m00 z   an vdd vdd p w=1.54u  l=0.13u ad=0.325998p pd=2.02012u as=0.35882p  ps=2.28709u
m01 vdd an z   vdd p w=1.54u  l=0.13u ad=0.35882p  pd=2.28709u as=0.325998p ps=2.02012u
m02 z   an vdd vdd p w=1.54u  l=0.13u ad=0.325998p pd=2.02012u as=0.35882p  ps=2.28709u
m03 vdd an z   vdd p w=1.54u  l=0.13u ad=0.35882p  pd=2.28709u as=0.325998p ps=2.02012u
m04 z   an vdd vdd p w=1.54u  l=0.13u ad=0.325998p pd=2.02012u as=0.35882p  ps=2.28709u
m05 vdd an z   vdd p w=1.265u l=0.13u ad=0.294745p pd=1.87868u as=0.267784p ps=1.65939u
m06 an  a  vdd vdd p w=1.045u l=0.13u ad=0.264825p pd=1.92333u as=0.243485p ps=1.55195u
m07 vdd a  an  vdd p w=1.045u l=0.13u ad=0.243485p pd=1.55195u as=0.264825p ps=1.92333u
m08 an  a  vdd vdd p w=1.045u l=0.13u ad=0.264825p pd=1.92333u as=0.243485p ps=1.55195u
m09 z   an vss vss n w=1.1u   l=0.13u ad=0.231p    pd=1.52u    as=0.304464p ps=2.08036u
m10 vss an z   vss n w=1.1u   l=0.13u ad=0.304464p pd=2.08036u as=0.231p    ps=1.52u   
m11 z   an vss vss n w=1.1u   l=0.13u ad=0.231p    pd=1.52u    as=0.304464p ps=2.08036u
m12 vss an z   vss n w=1.1u   l=0.13u ad=0.304464p pd=2.08036u as=0.231p    ps=1.52u   
m13 an  a  vss vss n w=0.88u  l=0.13u ad=0.1848p   pd=1.3u     as=0.243571p ps=1.66429u
m14 vss a  an  vss n w=0.88u  l=0.13u ad=0.243571p pd=1.66429u as=0.1848p   ps=1.3u    
C0 vdd an  0.129f
C1 vdd z   0.077f
C2 vdd a   0.008f
C3 an  z   0.242f
C4 an  a   0.167f
C5 a   vss 0.219f
C6 z   vss 0.322f
C7 an  vss 0.495f
.ends
