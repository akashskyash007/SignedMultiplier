.subckt cgi2v0x2 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from cgi2v0x2.ext -        technology: scmos
m00 n1  a vdd vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.464567p  ps=2.65667u 
m01 z   c n1  vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.3234p    ps=1.96u    
m02 n1  c z   vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.3234p    ps=1.96u    
m03 vdd a n1  vdd p w=1.54u  l=0.13u ad=0.464567p  pd=2.65667u as=0.3234p    ps=1.96u    
m04 w1  a vdd vdd p w=1.54u  l=0.13u ad=0.19635p   pd=1.795u   as=0.464567p  ps=2.65667u 
m05 z   b w1  vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.19635p   ps=1.795u   
m06 w2  b z   vdd p w=1.54u  l=0.13u ad=0.19635p   pd=1.795u   as=0.3234p    ps=1.96u    
m07 vdd a w2  vdd p w=1.54u  l=0.13u ad=0.464567p  pd=2.65667u as=0.19635p   ps=1.795u   
m08 n1  b vdd vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.464567p  ps=2.65667u 
m09 vdd b n1  vdd p w=1.54u  l=0.13u ad=0.464567p  pd=2.65667u as=0.3234p    ps=1.96u    
m10 n3  a vss vss n w=0.77u  l=0.13u ad=0.1617p    pd=1.19u    as=0.286733p  ps=1.96u    
m11 z   c n3  vss n w=0.77u  l=0.13u ad=0.166238p  pd=1.2725u  as=0.1617p    ps=1.19u    
m12 n3  c z   vss n w=0.77u  l=0.13u ad=0.1617p    pd=1.19u    as=0.166238p  ps=1.2725u  
m13 vss a n3  vss n w=0.77u  l=0.13u ad=0.286733p  pd=1.96u    as=0.1617p    ps=1.19u    
m14 w3  a vss vss n w=0.935u l=0.13u ad=0.119213p  pd=1.19u    as=0.348176p  ps=2.38u    
m15 z   b w3  vss n w=0.935u l=0.13u ad=0.20186p   pd=1.54518u as=0.119213p  ps=1.19u    
m16 w4  b z   vss n w=0.605u l=0.13u ad=0.0771375p pd=0.86u    as=0.130615p  ps=0.999821u
m17 vss a w4  vss n w=0.605u l=0.13u ad=0.225291p  pd=1.54u    as=0.0771375p ps=0.86u    
m18 n3  b vss vss n w=0.77u  l=0.13u ad=0.1617p    pd=1.19u    as=0.286733p  ps=1.96u    
m19 vss b n3  vss n w=0.77u  l=0.13u ad=0.286733p  pd=1.96u    as=0.1617p    ps=1.19u    
C0  a   n1  0.289f
C1  c   vdd 0.014f
C2  w4  n3  0.004f
C3  a   z   0.276f
C4  c   n1  0.022f
C5  b   vdd 0.028f
C6  w3  z   0.006f
C7  c   z   0.147f
C8  a   w1  0.009f
C9  b   n1  0.023f
C10 b   z   0.059f
C11 a   w2  0.015f
C12 vdd n1  0.302f
C13 a   n3  0.019f
C14 vdd z   0.017f
C15 w3  n3  0.008f
C16 c   n3  0.012f
C17 n1  z   0.046f
C18 vdd w1  0.004f
C19 w4  b   0.007f
C20 b   n3  0.099f
C21 n1  w1  0.008f
C22 vdd w2  0.004f
C23 z   w1  0.006f
C24 n1  w2  0.008f
C25 a   c   0.263f
C26 a   b   0.414f
C27 z   n3  0.191f
C28 a   vdd 0.125f
C29 w4  vss 0.002f
C30 w3  vss 0.004f
C31 n3  vss 0.426f
C32 w2  vss 0.006f
C33 w1  vss 0.007f
C34 z   vss 0.131f
C35 n1  vss 0.071f
C37 b   vss 0.295f
C38 c   vss 0.142f
C39 a   vss 0.425f
.ends
