.subckt vddtie vdd vss z
*10-JAN-08 SPICE3       file   created      from vddtie.ext -        technology: scmos
m00 z   vss vdd vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 vdd vss z   vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 z   vss w1  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m03 w2  vss z   vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0 vdd z   0.054f
C1 w2  vss 0.014f
C2 w1  vss 0.014f
C3 z   vss 0.115f
.ends
