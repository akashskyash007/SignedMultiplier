.subckt vfeed5 vdd vss
*01-JAN-08 SPICE3       file   created      from vfeed5.ext -        technology: scmos
.ends
