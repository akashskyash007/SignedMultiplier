.subckt vfeed5 vdd vss
*04-JAN-08 SPICE3       file   created      from vfeed5.ext -        technology: scmos
.ends
