.subckt nd2av0x05 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2av0x05.ext -        technology: scmos
m00 z   b  vdd vdd p w=0.44u  l=0.13u ad=0.0924p    pd=0.86u    as=0.287862p  ps=2.31692u
m01 vdd an z   vdd p w=0.44u  l=0.13u ad=0.287862p  pd=2.31692u as=0.0924p    ps=0.86u   
m02 an  a  vdd vdd p w=0.55u  l=0.13u ad=0.18205p   pd=1.85u    as=0.359827p  ps=2.89615u
m03 w1  b  z   vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u    as=0.144375p  ps=1.52u   
m04 vss an w1  vss n w=0.385u l=0.13u ad=0.263281p  pd=1.93308u as=0.0490875p ps=0.64u   
m05 an  a  vss vss n w=0.33u  l=0.13u ad=0.12375p   pd=1.41u    as=0.225669p  ps=1.65692u
C0  b   z   0.067f
C1  a   an  0.191f
C2  a   z   0.007f
C3  an  z   0.104f
C4  z   w1  0.007f
C5  vdd b   0.092f
C6  vdd an  0.014f
C7  vdd z   0.008f
C8  b   an  0.063f
C9  z   vss 0.053f
C10 an  vss 0.219f
C11 a   vss 0.115f
C12 b   vss 0.142f
.ends
