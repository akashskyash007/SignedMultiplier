.subckt nd2av0x2 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from nd2av0x2.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.54u l=0.13u ad=0.54725p  pd=3.28u as=0.5775p   ps=3.83u
m01 w2  a   vdd vdd p w=1.54u l=0.13u ad=0.5775p   pd=3.83u as=0.54725p  ps=3.28u
m02 z   w2  vdd vdd p w=1.54u l=0.13u ad=0.517p    pd=2.73u as=0.54725p  ps=3.28u
m03 vdd b   z   vdd p w=1.54u l=0.13u ad=0.54725p  pd=3.28u as=0.517p    ps=2.73u
m04 vss vdd w3  vss n w=1.1u  l=0.13u ad=0.404433p pd=2.51u as=0.4125p   ps=2.95u
m05 w2  a   vss vss n w=1.1u  l=0.13u ad=0.4125p   pd=2.95u as=0.404433p ps=2.51u
m06 w4  w2  vss vss n w=1.1u  l=0.13u ad=0.4004p   pd=2.29u as=0.404433p ps=2.51u
m07 z   b   w4  vss n w=1.1u  l=0.13u ad=0.4125p   pd=2.95u as=0.4004p   ps=2.29u
C0  w2  z   0.047f
C1  w2  b   0.089f
C2  z   b   0.126f
C3  z   w4  0.022f
C4  vdd a   0.130f
C5  vdd w2  0.038f
C6  vdd z   0.018f
C7  vdd b   0.038f
C8  a   w2  0.075f
C9  w4  vss 0.023f
C10 w3  vss 0.014f
C11 w1  vss 0.019f
C12 b   vss 0.153f
C13 z   vss 0.084f
C14 w2  vss 0.272f
C15 a   vss 0.179f
.ends
