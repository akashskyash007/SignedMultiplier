.subckt nd2v0x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v0x1.ext -        technology: scmos
m00 z   b vdd vdd p w=0.77u l=0.13u ad=0.1617p  pd=1.19u  as=0.34925p ps=2.51u 
m01 vdd a z   vdd p w=0.77u l=0.13u ad=0.34925p pd=2.51u  as=0.1617p  ps=1.19u 
m02 w1  b z   vss n w=0.66u l=0.13u ad=0.08415p pd=0.915u as=0.2112p  ps=2.07u 
m03 vss a w1  vss n w=0.66u l=0.13u ad=0.429p   pd=2.62u  as=0.08415p ps=0.915u
C0 vdd z   0.080f
C1 b   a   0.119f
C2 b   z   0.071f
C3 a   z   0.008f
C4 w1  vss 0.008f
C5 z   vss 0.186f
C6 a   vss 0.142f
C7 b   vss 0.113f
.ends
