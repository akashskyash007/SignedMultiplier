.subckt noa2a22_x1 i0 i1 i2 i3 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa2a22_x1.ext -        technology: scmos
m00 nq  i0 w1  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.728325p ps=3.975u
m01 w1  i1 nq  vdd p w=2.19u l=0.13u ad=0.728325p pd=3.975u as=0.58035p  ps=2.72u 
m02 vdd i3 w1  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.728325p ps=3.975u
m03 w1  i2 vdd vdd p w=2.19u l=0.13u ad=0.728325p pd=3.975u as=0.58035p  ps=2.72u 
m04 w2  i0 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u  as=0.46325p  ps=3.03u 
m05 nq  i1 w2  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u  as=0.28885p  ps=1.62u 
m06 w3  i3 nq  vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u  as=0.28885p  ps=1.62u 
m07 vss i2 w3  vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u  as=0.28885p  ps=1.62u 
C0  i1  w1  0.005f
C1  i3  i2  0.247f
C2  i1  nq  0.146f
C3  i3  w1  0.014f
C4  i3  nq  0.140f
C5  i2  w1  0.034f
C6  vdd i0  0.010f
C7  i1  w2  0.015f
C8  w1  nq  0.087f
C9  vdd i1  0.010f
C10 vdd i3  0.044f
C11 i3  w3  0.015f
C12 vdd i2  0.035f
C13 i0  i1  0.221f
C14 vdd w1  0.193f
C15 vdd nq  0.019f
C16 i1  i3  0.096f
C17 i0  w1  0.014f
C18 w3  vss 0.027f
C19 w2  vss 0.027f
C20 nq  vss 0.128f
C21 w1  vss 0.084f
C22 i2  vss 0.162f
C23 i3  vss 0.159f
C24 i1  vss 0.154f
C25 i0  vss 0.158f
.ends
