.subckt xoon21v0x1 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from xoon21v0x1.ext -        technology: scmos
m00 z   an bn  vdd p w=1.54u  l=0.13u ad=0.3234p    pd=1.96u    as=0.4444p    ps=3.83u   
m01 an  bn z   vdd p w=1.54u  l=0.13u ad=0.3619p    pd=2.57818u as=0.3234p    ps=1.96u   
m02 w1  a2 an  vdd p w=1.485u l=0.13u ad=0.189338p  pd=1.74u    as=0.348975p  ps=2.4861u 
m03 vdd a1 w1  vdd p w=1.485u l=0.13u ad=0.473079p  pd=2.79468u as=0.189338p  ps=1.74u   
m04 w2  a2 an  vdd p w=1.21u  l=0.13u ad=0.154275p  pd=1.465u   as=0.28435p   ps=2.02571u
m05 vdd a1 w2  vdd p w=1.21u  l=0.13u ad=0.385471p  pd=2.27714u as=0.154275p  ps=1.465u  
m06 bn  b  vdd vdd p w=1.54u  l=0.13u ad=0.4444p    pd=3.83u    as=0.4906p    ps=2.89818u
m07 w3  an vss vss n w=0.715u l=0.13u ad=0.0911625p pd=0.97u    as=0.256559p  ps=1.85824u
m08 z   bn w3  vss n w=0.715u l=0.13u ad=0.15015p   pd=1.135u   as=0.0911625p ps=0.97u   
m09 an  b  z   vss n w=0.715u l=0.13u ad=0.199824p  pd=1.67289u as=0.15015p   ps=1.135u  
m10 vss a2 an  vss n w=0.66u  l=0.13u ad=0.236824p  pd=1.71529u as=0.184453p  ps=1.54421u
m11 vss a1 an  vss n w=0.715u l=0.13u ad=0.256559p  pd=1.85824u as=0.199824p  ps=1.67289u
m12 bn  b  vss vss n w=0.715u l=0.13u ad=0.225775p  pd=2.18u    as=0.256559p  ps=1.85824u
C0  an  z   0.204f
C1  vdd a1  0.036f
C2  an  a2  0.100f
C3  bn  z   0.082f
C4  vdd w1  0.003f
C5  an  a1  0.011f
C6  vdd b   0.036f
C7  bn  a2  0.099f
C8  bn  a1  0.038f
C9  an  b   0.004f
C10 bn  w1  0.036f
C11 bn  b   0.155f
C12 a2  a1  0.209f
C13 bn  w2  0.008f
C14 vdd an  0.019f
C15 a2  b   0.041f
C16 vdd bn  0.281f
C17 z   w3  0.009f
C18 a2  w2  0.019f
C19 a1  b   0.126f
C20 vdd z   0.007f
C21 vdd a2  0.009f
C22 an  bn  0.350f
C23 w3  vss 0.007f
C24 w2  vss 0.003f
C25 b   vss 0.235f
C26 w1  vss 0.004f
C27 a1  vss 0.183f
C28 a2  vss 0.168f
C29 z   vss 0.255f
C30 bn  vss 0.312f
C31 an  vss 0.288f
.ends
