.subckt or3v0x05 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from or3v0x05.ext -        technology: scmos
m00 vdd zn z   vdd p w=0.66u  l=0.13u ad=0.188635p pd=1.2u    as=0.2112p   ps=2.07u  
m01 w1  a  vdd vdd p w=1.375u l=0.13u ad=0.175313p pd=1.63u   as=0.39299p  ps=2.5u   
m02 w2  b  w1  vdd p w=1.375u l=0.13u ad=0.175313p pd=1.63u   as=0.175313p ps=1.63u  
m03 zn  c  w2  vdd p w=1.375u l=0.13u ad=0.400675p pd=3.5u    as=0.175313p ps=1.63u  
m04 vss zn z   vss n w=0.33u  l=0.13u ad=0.119213p pd=1.0525u as=0.12375p  ps=1.41u  
m05 zn  a  vss vss n w=0.33u  l=0.13u ad=0.08745p  pd=0.97u   as=0.119213p ps=1.0525u
m06 vss b  zn  vss n w=0.33u  l=0.13u ad=0.119213p pd=1.0525u as=0.08745p  ps=0.97u  
m07 zn  c  vss vss n w=0.33u  l=0.13u ad=0.08745p  pd=0.97u   as=0.119213p ps=1.0525u
C0  vdd z   0.034f
C1  a   c   0.029f
C2  vdd w1  0.003f
C3  a   zn  0.154f
C4  b   c   0.152f
C5  a   z   0.007f
C6  b   zn  0.072f
C7  vdd w2  0.003f
C8  a   w1  0.006f
C9  c   zn  0.085f
C10 zn  z   0.111f
C11 c   w2  0.012f
C12 zn  w1  0.022f
C13 vdd a   0.007f
C14 zn  w2  0.008f
C15 vdd b   0.007f
C16 vdd c   0.007f
C17 vdd zn  0.094f
C18 a   b   0.131f
C19 w2  vss 0.007f
C20 w1  vss 0.006f
C21 z   vss 0.213f
C22 zn  vss 0.322f
C23 c   vss 0.117f
C24 b   vss 0.108f
C25 a   vss 0.108f
.ends
