.subckt an2v2x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from an2v2x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.423127p pd=2.95355u as=0.48675p  ps=3.83u   
m01 zn  a  vdd vdd p w=0.935u l=0.13u ad=0.19635p  pd=1.355u   as=0.256899p ps=1.79323u
m02 vdd b  zn  vdd p w=0.935u l=0.13u ad=0.256899p pd=1.79323u as=0.19635p  ps=1.355u  
m03 vss zn z   vss n w=0.77u  l=0.13u ad=0.320513p pd=1.85u    as=0.28875p  ps=2.29u   
m04 w1  a  vss vss n w=0.77u  l=0.13u ad=0.098175p pd=1.025u   as=0.320513p ps=1.85u   
m05 zn  b  w1  vss n w=0.77u  l=0.13u ad=0.24035p  pd=2.29u    as=0.098175p ps=1.025u  
C0  vdd a   0.006f
C1  vdd b   0.021f
C2  zn  w1  0.008f
C3  a   b   0.151f
C4  a   w1  0.007f
C5  zn  z   0.158f
C6  zn  vdd 0.052f
C7  zn  a   0.148f
C8  z   vdd 0.024f
C9  zn  b   0.028f
C10 z   a   0.006f
C11 w1  vss 0.003f
C12 b   vss 0.095f
C13 a   vss 0.099f
C15 z   vss 0.228f
C16 zn  vss 0.225f
.ends
