.subckt no2_x1 i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from no2_x1.ext -        technology: scmos
m00 w1  i1 nq  vdd p w=2.09u l=0.13u ad=0.32395p pd=2.4u  as=1.18608p ps=5.59u
m01 vdd i0 w1  vdd p w=2.09u l=0.13u ad=0.8987p  pd=5.04u as=0.32395p ps=2.4u 
m02 nq  i1 vss vss n w=0.55u l=0.13u ad=0.14575p pd=1.08u as=0.3817p  ps=2.84u
m03 vss i0 nq  vss n w=0.55u l=0.13u ad=0.3817p  pd=2.84u as=0.14575p ps=1.08u
C0  i1 i0  0.273f
C1  i1 nq  0.183f
C2  i0 nq  0.012f
C3  i1 w1  0.019f
C4  i1 vdd 0.023f
C5  i0 vdd 0.054f
C6  nq vdd 0.021f
C7  w1 vdd 0.010f
C9  w1 vss 0.011f
C10 nq vss 0.176f
C11 i0 vss 0.189f
C12 i1 vss 0.141f
.ends
