* Spice description of vddtie
* Spice driver version 134999461
* Date  4/01/2008 at 19:50:04
* vsxlib 0.13um values
.subckt vddtie vdd vss z
M1  z     vss   vdd   vdd p  L=0.12U  W=1.65U  AS=0.43725P  AD=0.43725P  PS=3.83U   PD=3.83U
M2  vss   vss   z     vss n  L=0.12U  W=1.265U AS=0.335225P AD=0.335225P PS=3.06U   PD=3.06U
C1  z     vss   0.828f
.ends
