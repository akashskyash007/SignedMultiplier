* Spice description of oan21_x2
* Spice driver version 134999461
* Date  4/01/2008 at 19:11:41
* vxlib 0.13um values
.subckt oan21_x2 a1 a2 b vdd vss z
M1  n1    a1    vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2_1 z     sig1  vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2  sig1  a2    n1    vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M3  vdd   b     sig1  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M4  n2    a1    vss   vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M5  vss   a2    n2    vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M6_2 z     sig1  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M6  n2    b     sig1  vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
C7  a1    vss   0.836f
C8  a2    vss   0.814f
C9  b     vss   0.842f
C2  n2    vss   0.262f
C1  sig1  vss   0.976f
C4  z     vss   0.673f
.ends
