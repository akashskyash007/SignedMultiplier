* Spice description of iv1_w2
* Spice driver version 134999461
* Date  4/01/2008 at 18:59:12
* vxlib 0.13um values
.subckt iv1_w2 a vdd vss z
M1  vdd   a     z     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
M2  z     a     vss   vss n  L=0.12U  W=1.43U  AS=0.37895P  AD=0.37895P  PS=3.39U   PD=3.39U
C4  a     vss   0.561f
C2  z     vss   0.618f
.ends
