.subckt cgi2abv0x05 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from cgi2abv0x05.ext -        technology: scmos
m00 vdd a  an  vdd p w=1.1u   l=0.13u ad=0.275p     pd=1.95227u as=0.37015p   ps=2.95u   
m01 n1  an vdd vdd p w=0.88u  l=0.13u ad=0.22715p   pd=1.70333u as=0.22p      ps=1.56182u
m02 w1  an vdd vdd p w=0.88u  l=0.13u ad=0.1122p    pd=1.135u   as=0.22p      ps=1.56182u
m03 z   bn w1  vdd p w=0.88u  l=0.13u ad=0.1848p    pd=1.3u     as=0.1122p    ps=1.135u  
m04 n1  c  z   vdd p w=0.88u  l=0.13u ad=0.22715p   pd=1.70333u as=0.1848p    ps=1.3u    
m05 vdd bn n1  vdd p w=0.88u  l=0.13u ad=0.22p      pd=1.56182u as=0.22715p   ps=1.70333u
m06 bn  b  vdd vdd p w=1.1u   l=0.13u ad=0.37015p   pd=2.95u    as=0.275p     ps=1.95227u
m07 vss a  an  vss n w=0.55u  l=0.13u ad=0.251994p  pd=2.09512u as=0.18205p   ps=1.85u   
m08 w2  an vss vss n w=0.385u l=0.13u ad=0.0490875p pd=0.64u    as=0.176396p  ps=1.46659u
m09 z   bn w2  vss n w=0.385u l=0.13u ad=0.08085p   pd=0.805u   as=0.0490875p ps=0.64u   
m10 n3  c  z   vss n w=0.385u l=0.13u ad=0.102025p  pd=1.04333u as=0.08085p   ps=0.805u  
m11 vss bn n3  vss n w=0.385u l=0.13u ad=0.176396p  pd=1.46659u as=0.102025p  ps=1.04333u
m12 n3  an vss vss n w=0.385u l=0.13u ad=0.102025p  pd=1.04333u as=0.176396p  ps=1.46659u
m13 bn  b  vss vss n w=0.55u  l=0.13u ad=0.18205p   pd=1.85u    as=0.251994p  ps=2.09512u
C0  w1  z   0.002f
C1  vdd n1  0.142f
C2  an  bn  0.106f
C3  z   w2  0.008f
C4  bn  c   0.223f
C5  z   n3  0.062f
C6  an  n1  0.017f
C7  bn  b   0.185f
C8  bn  n1  0.006f
C9  an  z   0.025f
C10 c   n1  0.038f
C11 bn  z   0.020f
C12 vdd an  0.070f
C13 c   z   0.109f
C14 an  n3  0.005f
C15 vdd bn  0.061f
C16 bn  n3  0.020f
C17 n1  w1  0.022f
C18 vdd c   0.002f
C19 a   an  0.183f
C20 c   n3  0.007f
C21 n1  z   0.073f
C22 vdd b   0.008f
C23 n3  vss 0.236f
C24 z   vss 0.057f
C25 w1  vss 0.003f
C26 n1  vss 0.047f
C27 b   vss 0.109f
C28 c   vss 0.113f
C29 bn  vss 0.254f
C30 an  vss 0.307f
C31 a   vss 0.135f
.ends
