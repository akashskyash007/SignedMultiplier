* Spice description of iv1v4x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:45:37
* vsclib 0.13um values
.subckt iv1v4x2 a vdd vss z
M01 z     a     vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 vdd   a     z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M03 vss   a     z     vss n  L=0.12U  W=0.44U  AS=0.1166P   AD=0.1166P   PS=1.41U   PD=1.41U
C3  a     vss   0.546f
C1  z     vss   0.448f
.ends
