* Spice description of vfeed2
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:39
* wsclib 0.13um values
.subckt vfeed2 vdd vss
.ends
