.subckt oan21v0x05 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from oan21v0x05.ext -        technology: scmos
m00 vdd zn z   vdd p w=0.66u  l=0.13u ad=0.478783p  pd=2.35543u  as=0.2112p   ps=2.07u   
m01 zn  b  vdd vdd p w=0.44u  l=0.13u ad=0.0997652p pd=0.866087u as=0.319189p ps=1.57029u
m02 w1  a2 zn  vdd p w=0.825u l=0.13u ad=0.105188p  pd=1.08u     as=0.18706p  ps=1.62391u
m03 vdd a1 w1  vdd p w=0.825u l=0.13u ad=0.598479p  pd=2.94429u  as=0.105188p ps=1.08u   
m04 vss zn z   vss n w=0.33u  l=0.13u ad=0.18546p   pd=1.5u      as=0.12375p  ps=1.41u   
m05 n1  b  zn  vss n w=0.385u l=0.13u ad=0.102025p  pd=1.04333u  as=0.144375p ps=1.52u   
m06 vss a2 n1  vss n w=0.385u l=0.13u ad=0.21637p   pd=1.75u     as=0.102025p ps=1.04333u
m07 n1  a1 vss vss n w=0.385u l=0.13u ad=0.102025p  pd=1.04333u  as=0.21637p  ps=1.75u   
C0  vdd z   0.015f
C1  a2  b   0.081f
C2  vdd w1  0.003f
C3  a1  b   0.014f
C4  b   zn  0.061f
C5  a2  n1  0.059f
C6  a1  n1  0.006f
C7  b   w1  0.003f
C8  zn  z   0.035f
C9  vdd a2  0.007f
C10 zn  n1  0.011f
C11 vdd a1  0.013f
C12 vdd zn  0.103f
C13 a2  a1  0.104f
C14 n1  vss 0.148f
C15 w1  vss 0.005f
C16 z   vss 0.160f
C17 zn  vss 0.148f
C18 b   vss 0.109f
C19 a1  vss 0.124f
C20 a2  vss 0.114f
.ends
