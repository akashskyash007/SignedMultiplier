.subckt cgi2v0x3 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from cgi2v0x3.ext -        technology: scmos
m00 n1  b vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u as=0.398689p ps=2.22889u
m01 vdd b n1  vdd p w=1.54u l=0.13u ad=0.398689p pd=2.22889u as=0.34155p  ps=2.16778u
m02 n1  b vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u as=0.398689p ps=2.22889u
m03 z   c n1  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u    as=0.34155p  ps=2.16778u
m04 n1  c z   vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u as=0.3234p   ps=1.96u   
m05 z   c n1  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u    as=0.34155p  ps=2.16778u
m06 w1  b z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m07 vdd a w1  vdd p w=1.54u l=0.13u ad=0.398689p pd=2.22889u as=0.19635p  ps=1.795u  
m08 w2  a vdd vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.398689p ps=2.22889u
m09 z   b w2  vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u    as=0.19635p  ps=1.795u  
m10 w3  b z   vdd p w=1.54u l=0.13u ad=0.19635p  pd=1.795u   as=0.3234p   ps=1.96u   
m11 vdd a w3  vdd p w=1.54u l=0.13u ad=0.398689p pd=2.22889u as=0.19635p  ps=1.795u  
m12 n1  a vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u as=0.398689p ps=2.22889u
m13 vdd a n1  vdd p w=1.54u l=0.13u ad=0.398689p pd=2.22889u as=0.34155p  ps=2.16778u
m14 n1  a vdd vdd p w=1.54u l=0.13u ad=0.34155p  pd=2.16778u as=0.398689p ps=2.22889u
m15 n3  b vss vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u as=0.263818p ps=1.67097u
m16 vss b n3  vss n w=0.77u l=0.13u ad=0.263818p pd=1.67097u as=0.1617p   ps=1.14935u
m17 n3  b vss vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u as=0.263818p ps=1.67097u
m18 z   c n3  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u    as=0.1617p   ps=1.14935u
m19 n3  c z   vss n w=0.77u l=0.13u ad=0.1617p   pd=1.14935u as=0.1617p   ps=1.19u   
m20 z   c n3  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u    as=0.1617p   ps=1.14935u
m21 w4  b z   vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u   as=0.1617p   ps=1.19u   
m22 vss a w4  vss n w=0.77u l=0.13u ad=0.263818p pd=1.67097u as=0.098175p ps=1.025u  
m23 w5  a vss vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u   as=0.263818p ps=1.67097u
m24 z   b w5  vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u    as=0.098175p ps=1.025u  
m25 w6  b z   vss n w=0.77u l=0.13u ad=0.098175p pd=1.025u   as=0.1617p   ps=1.19u   
m26 vss a w6  vss n w=0.77u l=0.13u ad=0.263818p pd=1.67097u as=0.098175p ps=1.025u  
m27 n3  a vss vss n w=1.1u  l=0.13u ad=0.231p    pd=1.64194u as=0.376883p ps=2.3871u 
m28 vss a n3  vss n w=1.1u  l=0.13u ad=0.376883p pd=2.3871u  as=0.231p    ps=1.64194u
C0  a   z   0.291f
C1  n3  b   0.119f
C2  n1  z   0.388f
C3  n3  c   0.036f
C4  a   w2  0.006f
C5  n1  w1  0.008f
C6  vdd b   0.042f
C7  n3  a   0.030f
C8  a   w3  0.006f
C9  z   w1  0.009f
C10 n1  w2  0.008f
C11 vdd c   0.021f
C12 n3  w4  0.008f
C13 z   w2  0.009f
C14 n1  w3  0.008f
C15 vdd a   0.061f
C16 n3  z   0.337f
C17 w6  z   0.009f
C18 z   w3  0.009f
C19 vdd n1  0.480f
C20 b   c   0.204f
C21 vdd z   0.081f
C22 b   a   0.553f
C23 n3  w5  0.008f
C24 b   n1  0.031f
C25 vdd w1  0.004f
C26 n3  w6  0.008f
C27 w4  b   0.006f
C28 b   z   0.078f
C29 c   n1  0.023f
C30 vdd w2  0.004f
C31 c   z   0.155f
C32 a   n1  0.037f
C33 vdd w3  0.004f
C34 w5  b   0.007f
C35 w6  vss 0.003f
C36 w5  vss 0.004f
C37 w4  vss 0.004f
C38 n3  vss 0.538f
C39 w3  vss 0.006f
C40 w2  vss 0.007f
C41 w1  vss 0.007f
C42 z   vss 0.220f
C43 n1  vss 0.154f
C44 a   vss 0.386f
C45 c   vss 0.194f
C46 b   vss 0.522f
.ends
