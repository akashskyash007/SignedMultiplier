.subckt a4_x4 i0 i1 i2 i3 q vdd vss
*05-JAN-08 SPICE3       file   created      from a4_x4.ext -        technology: scmos
m00 w1  i0 vdd vdd p w=1.1u   l=0.13u ad=0.293827p pd=1.6718u  as=0.388143p ps=2.47013u
m01 vdd i1 w1  vdd p w=1.1u   l=0.13u ad=0.388143p pd=2.47013u as=0.293827p ps=1.6718u 
m02 w1  i2 vdd vdd p w=1.045u l=0.13u ad=0.279136p pd=1.58821u as=0.368736p ps=2.34662u
m03 vdd i3 w1  vdd p w=1.045u l=0.13u ad=0.368736p pd=2.34662u as=0.279136p ps=1.58821u
m04 q   w1 vdd vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.737471p ps=4.69325u
m05 vdd w1 q   vdd p w=2.09u  l=0.13u ad=0.737471p pd=4.69325u as=0.55385p  ps=2.62u   
m06 w2  i0 vss vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.46145p  ps=3.28u   
m07 w3  i1 w2  vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.161975p ps=1.355u  
m08 w4  i2 w3  vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.161975p ps=1.355u  
m09 w1  i3 w4  vss n w=1.045u l=0.13u ad=0.36465p  pd=2.95u    as=0.161975p ps=1.355u  
m10 q   w1 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.46145p  ps=3.28u   
m11 vss w1 q   vss n w=1.045u l=0.13u ad=0.46145p  pd=3.28u    as=0.276925p ps=1.575u  
C0  i2  i3  0.223f
C1  i1  w2  0.012f
C2  i1  w3  0.012f
C3  vdd w1  0.188f
C4  vdd i0  0.013f
C5  i2  w4  0.020f
C6  vdd i1  0.004f
C7  w1  i1  0.035f
C8  vdd i2  0.018f
C9  w1  i2  0.028f
C10 vdd i3  0.003f
C11 i0  i1  0.264f
C12 vdd q   0.086f
C13 w1  i3  0.216f
C14 w1  q   0.219f
C15 i1  i2  0.266f
C16 w4  vss 0.005f
C17 w3  vss 0.006f
C18 w2  vss 0.006f
C19 q   vss 0.146f
C20 i3  vss 0.136f
C21 i2  vss 0.157f
C22 i1  vss 0.148f
C23 i0  vss 0.175f
C24 w1  vss 0.406f
.ends
