.subckt or3v0x4 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from or3v0x4.ext -        technology: scmos
m00 z   zn vdd vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.431922p ps=2.60094u
m01 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.431922p pd=2.60094u as=0.3234p   ps=1.96u   
m02 w1  a  vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.431922p ps=2.60094u
m03 w2  b  w1  vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.19635p  ps=1.795u  
m04 zn  c  w2  vdd p w=1.54u  l=0.13u ad=0.372808p pd=2.50056u as=0.19635p  ps=1.795u  
m05 w3  c  zn  vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.372808p ps=2.50056u
m06 w4  b  w3  vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.19635p  ps=1.795u  
m07 vdd a  w4  vdd p w=1.54u  l=0.13u ad=0.431922p pd=2.60094u as=0.19635p  ps=1.795u  
m08 w5  a  vdd vdd p w=0.88u  l=0.13u ad=0.1122p   pd=1.135u   as=0.246813p ps=1.48625u
m09 w6  b  w5  vdd p w=0.88u  l=0.13u ad=0.1122p   pd=1.135u   as=0.1122p   ps=1.135u  
m10 zn  c  w6  vdd p w=0.88u  l=0.13u ad=0.213033p pd=1.42889u as=0.1122p   ps=1.135u  
m11 z   zn vss vss n w=0.77u  l=0.13u ad=0.1617p   pd=1.19u    as=0.233758p ps=1.70299u
m12 vss zn z   vss n w=0.77u  l=0.13u ad=0.233758p pd=1.70299u as=0.1617p   ps=1.19u   
m13 zn  a  vss vss n w=0.715u l=0.13u ad=0.175358p pd=1.48333u as=0.217061p ps=1.58134u
m14 vss b  zn  vss n w=0.715u l=0.13u ad=0.217061p pd=1.58134u as=0.175358p ps=1.48333u
m15 zn  c  vss vss n w=0.715u l=0.13u ad=0.175358p pd=1.48333u as=0.217061p ps=1.58134u
C0  zn  w4  0.015f
C1  vdd zn  0.106f
C2  vdd a   0.014f
C3  vdd b   0.014f
C4  vdd c   0.014f
C5  zn  a   0.290f
C6  zn  b   0.099f
C7  vdd z   0.046f
C8  zn  c   0.071f
C9  vdd w1  0.004f
C10 a   b   0.398f
C11 zn  z   0.092f
C12 vdd w2  0.004f
C13 a   c   0.118f
C14 w6  zn  0.008f
C15 zn  w1  0.008f
C16 vdd w3  0.004f
C17 b   c   0.305f
C18 a   w1  0.006f
C19 zn  w2  0.008f
C20 vdd w4  0.004f
C21 a   w2  0.006f
C22 zn  w3  0.008f
C23 w5  zn  0.008f
C24 w6  vss 0.005f
C25 w5  vss 0.007f
C26 w4  vss 0.009f
C27 w3  vss 0.009f
C28 w2  vss 0.008f
C29 w1  vss 0.010f
C30 z   vss 0.214f
C31 c   vss 0.305f
C32 b   vss 0.256f
C33 a   vss 0.220f
C34 zn  vss 0.446f
.ends
