.subckt zero_x0 nq vdd vss
*05-JAN-08 SPICE3       file   created      from zero_x0.ext -        technology: scmos
m00 nq vdd vss vss n w=0.54u l=0.13u ad=0.2295p pd=1.93u as=0.2889p ps=2.15u
C0 vdd nq  0.124f
C1 nq  vss 0.137f
.ends
