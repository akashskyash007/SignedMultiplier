.subckt oa2a2a2a24_x4 i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss
*05-JAN-08 SPICE3       file   created      from oa2a2a2a24_x4.ext -        technology: scmos
m00 w1  i7 w2  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.75555p  ps=3.975u
m01 w2  i6 w1  vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.58035p  ps=2.72u 
m02 w2  i5 w3  vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.75555p  ps=3.975u
m03 w3  i4 w2  vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.75555p  ps=3.975u
m04 w4  i3 w3  vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.75555p  ps=3.975u
m05 w3  i2 w4  vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.58035p  ps=2.72u 
m06 w4  i1 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.75555p  ps=3.975u
m07 vdd i0 w4  vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.58035p  ps=2.72u 
m08 q   w1 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u  as=0.75555p  ps=3.975u
m09 vdd w1 q   vdd p w=2.19u l=0.13u ad=0.75555p  pd=3.975u as=0.58035p  ps=2.72u 
m10 w5  i7 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u  as=0.405117p ps=2.56u 
m11 w1  i6 w5  vss n w=1.09u l=0.13u ad=0.37605p  pd=2.325u as=0.28885p  ps=1.62u 
m12 w6  i5 vss vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u   as=0.405117p ps=2.56u 
m13 w1  i4 w6  vss n w=1.09u l=0.13u ad=0.37605p  pd=2.325u as=0.16895p  ps=1.4u  
m14 w7  i3 w1  vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u   as=0.37605p  ps=2.325u
m15 vss i2 w7  vss n w=1.09u l=0.13u ad=0.405117p pd=2.56u  as=0.16895p  ps=1.4u  
m16 w8  i1 w1  vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u   as=0.37605p  ps=2.325u
m17 vss i0 w8  vss n w=1.09u l=0.13u ad=0.405117p pd=2.56u  as=0.16895p  ps=1.4u  
m18 q   w1 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u  as=0.405117p ps=2.56u 
m19 vss w1 q   vss n w=1.09u l=0.13u ad=0.405117p pd=2.56u  as=0.28885p  ps=1.62u 
C0  w1  i7  0.095f
C1  w1  w6  0.008f
C2  w4  vdd 0.084f
C3  i1  i0  0.113f
C4  w1  i6  0.091f
C5  w2  i7  0.014f
C6  i5  i4  0.227f
C7  w1  w7  0.008f
C8  i1  w1  0.060f
C9  w1  i5  0.014f
C10 w2  i6  0.030f
C11 i2  w1  0.019f
C12 vdd q   0.070f
C13 i0  w1  0.121f
C14 w1  i4  0.014f
C15 w2  i5  0.023f
C16 i3  i2  0.227f
C17 w2  i4  0.005f
C18 w3  i5  0.005f
C19 vdd i7  0.010f
C20 i2  w3  0.005f
C21 i3  i4  0.195f
C22 i1  w4  0.014f
C23 w1  w2  0.041f
C24 w3  i4  0.010f
C25 vdd i6  0.010f
C26 i2  w4  0.029f
C27 i3  w1  0.014f
C28 i0  w4  0.005f
C29 i1  vdd 0.019f
C30 vdd i5  0.010f
C31 i2  vdd 0.010f
C32 w2  w3  0.074f
C33 i0  vdd 0.054f
C34 vdd i4  0.010f
C35 i7  i6  0.096f
C36 i3  w3  0.014f
C37 i0  q   0.114f
C38 w1  vdd 0.039f
C39 w1  q   0.007f
C40 w3  w4  0.066f
C41 w2  vdd 0.115f
C42 i3  vdd 0.010f
C43 w1  w5  0.011f
C44 w3  vdd 0.169f
C45 w8  vss 0.018f
C46 w7  vss 0.016f
C47 w6  vss 0.016f
C48 w5  vss 0.028f
C49 q   vss 0.137f
C51 w4  vss 0.060f
C52 w3  vss 0.089f
C53 w2  vss 0.108f
C54 w1  vss 0.707f
C55 i0  vss 0.131f
C56 i1  vss 0.123f
C57 i2  vss 0.122f
C58 i3  vss 0.130f
C59 i4  vss 0.118f
C60 i5  vss 0.129f
C61 i6  vss 0.142f
C62 i7  vss 0.157f
.ends
