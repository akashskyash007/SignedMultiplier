* Spice description of noa2a2a2a24_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:23:19
* ssxlib 0.13um values
.subckt noa2a2a2a24_x1 i0 i1 i2 i3 i4 i5 i6 i7 nq vdd vss
Mtr_00001 sig1  i7    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00002 sig12 i1    nq    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00003 sig6  i5    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00004 vss   i0    sig12 vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00005 vss   i2    sig9  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00006 nq    i6    sig1  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00007 sig9  i3    nq    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00008 nq    i4    sig6  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00009 sig15 i6    nq    vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00010 sig15 i5    sig16 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00011 sig16 i4    sig15 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00012 sig16 i2    sig17 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00013 vdd   i0    sig17 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00014 nq    i7    sig15 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00015 sig17 i1    vdd   vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
Mtr_00016 sig17 i3    sig16 vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
C14 i0    vss   0.726f
C13 i1    vss   0.726f
C10 i2    vss   0.685f
C11 i3    vss   0.628f
C8  i4    vss   0.628f
C7  i5    vss   0.628f
C5  i6    vss   0.703f
C4  i7    vss   0.726f
C2  nq    vss   1.209f
C15 sig15 vss   0.514f
C16 sig16 vss   0.401f
C17 sig17 vss   0.325f
.ends
