.subckt oai22_x05 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from oai22_x05.ext -        technology: scmos
m00 w1  b1 vdd vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u   as=0.6182p   ps=3.61u  
m01 z   b2 w1  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u   as=0.1705p   ps=1.41u  
m02 w2  a2 z   vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u   as=0.2915p   ps=1.63u  
m03 vdd a1 w2  vdd p w=1.1u   l=0.13u ad=0.6182p   pd=3.61u   as=0.1705p   ps=1.41u  
m04 z   b1 n3  vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u  as=0.1584p   ps=1.4375u
m05 n3  b2 z   vss n w=0.495u l=0.13u ad=0.1584p   pd=1.4375u as=0.131175p ps=1.025u 
m06 vss a2 n3  vss n w=0.495u l=0.13u ad=0.231p    pd=1.63u   as=0.1584p   ps=1.4375u
m07 n3  a1 vss vss n w=0.495u l=0.13u ad=0.1584p   pd=1.4375u as=0.231p    ps=1.63u  
C0  n3  w3  0.054f
C1  a1  z   0.023f
C2  b2  n3  0.046f
C3  vdd b1  0.004f
C4  w4  w3  0.166f
C5  vdd w3  0.043f
C6  b1  w5  0.010f
C7  a2  n3  0.022f
C8  a1  w2  0.024f
C9  w1  z   0.013f
C10 vdd b2  0.004f
C11 w5  w3  0.166f
C12 b2  w5  0.011f
C13 a2  w4  0.001f
C14 a1  n3  0.007f
C15 vdd a2  0.003f
C16 w6  w3  0.166f
C17 b1  w3  0.020f
C18 b2  w6  0.033f
C19 a2  w5  0.010f
C20 a1  w4  0.011f
C21 vdd a1  0.051f
C22 b1  b2  0.162f
C23 b2  w3  0.012f
C24 a2  w6  0.011f
C25 a1  w5  0.012f
C26 z   n3  0.046f
C27 a2  w3  0.017f
C28 a1  w6  0.001f
C29 z   w4  0.058f
C30 b1  a1  0.016f
C31 vdd z   0.115f
C32 b2  a2  0.168f
C33 a1  w3  0.017f
C34 z   w5  0.009f
C35 w2  w4  0.002f
C36 b1  w1  0.014f
C37 z   w6  0.030f
C38 b1  z   0.175f
C39 a2  a1  0.192f
C40 z   w3  0.025f
C41 vdd w4  0.013f
C42 b2  z   0.024f
C43 b1  n3  0.002f
C44 w3  vss 1.005f
C45 w6  vss 0.174f
C46 w5  vss 0.179f
C47 w4  vss 0.167f
C48 n3  vss 0.147f
C49 z   vss 0.043f
C50 a1  vss 0.071f
C51 a2  vss 0.092f
C52 b2  vss 0.099f
C53 b1  vss 0.082f
.ends
