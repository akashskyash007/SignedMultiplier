* Spice description of vfeed7
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:53
* vxlib 0.13um values
.subckt vfeed7 vdd vss
.ends
