.subckt bf1v8x4 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v8x4.ext -        technology: scmos
m00 z   an vdd vdd p w=1.54u l=0.13u ad=0.3234p   pd=1.96u    as=0.446921p ps=3.01389u
m01 vdd an z   vdd p w=1.54u l=0.13u ad=0.446921p pd=3.01389u as=0.3234p   ps=1.96u   
m02 an  a  vdd vdd p w=0.88u l=0.13u ad=0.31185p  pd=2.51u    as=0.255383p ps=1.72222u
m03 z   an vss vss n w=0.77u l=0.13u ad=0.1617p   pd=1.19u    as=0.206403p ps=1.81611u
m04 vss an z   vss n w=0.77u l=0.13u ad=0.206403p pd=1.81611u as=0.1617p   ps=1.19u   
m05 an  a  vss vss n w=0.44u l=0.13u ad=0.1529p   pd=1.63u    as=0.117944p ps=1.03778u
C0 vdd a   0.017f
C1 an  z   0.051f
C2 an  a   0.188f
C3 z   a   0.010f
C4 vdd an  0.045f
C5 vdd z   0.101f
C6 a   vss 0.087f
C7 z   vss 0.217f
C8 an  vss 0.252f
.ends
