.subckt nmx2_x4 cmd i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nmx2_x4.ext -        technology: scmos
m00 vdd cmd w1  vdd p w=1.09u l=0.13u ad=0.411369p pd=2.33215u as=0.46325p  ps=3.03u   
m01 w2  i0  vdd vdd p w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.411369p ps=2.33215u
m02 w3  cmd w2  vdd p w=1.09u l=0.13u ad=0.40875p  pd=1.84u    as=0.16895p  ps=1.4u    
m03 w4  w1  w3  vdd p w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.40875p  ps=1.84u   
m04 vdd i1  w4  vdd p w=1.09u l=0.13u ad=0.411369p pd=2.33215u as=0.16895p  ps=1.4u    
m05 w5  w3  vdd vdd p w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.411369p ps=2.33215u
m06 nq  w5  vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.826512p ps=4.6857u 
m07 vdd w5  nq  vdd p w=2.19u l=0.13u ad=0.826512p pd=4.6857u  as=0.58035p  ps=2.72u   
m08 vss cmd w1  vss n w=0.54u l=0.13u ad=0.186499p pd=1.28654u as=0.3703p   ps=2.81u   
m09 w6  i0  vss vss n w=0.54u l=0.13u ad=0.0837p   pd=0.85u    as=0.186499p ps=1.28654u
m10 w3  w1  w6  vss n w=0.54u l=0.13u ad=0.41535p  pd=2.28u    as=0.0837p   ps=0.85u   
m11 w7  cmd w3  vss n w=0.54u l=0.13u ad=0.0837p   pd=0.85u    as=0.41535p  ps=2.28u   
m12 vss i1  w7  vss n w=0.54u l=0.13u ad=0.186499p pd=1.28654u as=0.0837p   ps=0.85u   
m13 w5  w3  vss vss n w=0.54u l=0.13u ad=0.3703p   pd=2.81u    as=0.186499p ps=1.28654u
m14 nq  w5  vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.376452p ps=2.59691u
m15 vss w5  nq  vss n w=1.09u l=0.13u ad=0.376452p pd=2.59691u as=0.28885p  ps=1.62u   
C0  vdd i0  0.046f
C1  vdd w1  0.012f
C2  vdd i1  0.046f
C3  vdd w3  0.012f
C4  cmd i0  0.296f
C5  w5  i1  0.092f
C6  cmd w1  0.046f
C7  cmd i1  0.052f
C8  i0  w1  0.134f
C9  w5  w3  0.017f
C10 vdd nq  0.123f
C11 cmd w3  0.181f
C12 cmd w2  0.020f
C13 w1  i1  0.136f
C14 w5  nq  0.007f
C15 w1  w3  0.101f
C16 vdd w5  0.066f
C17 i1  w3  0.103f
C18 vdd cmd 0.015f
C19 w7  vss 0.012f
C20 w6  vss 0.012f
C21 nq  vss 0.136f
C22 w4  vss 0.010f
C23 w2  vss 0.006f
C24 w3  vss 0.254f
C25 i1  vss 0.179f
C26 w1  vss 0.440f
C27 i0  vss 0.152f
C28 cmd vss 0.339f
C29 w5  vss 0.299f
.ends
