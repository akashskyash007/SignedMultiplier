.subckt nr2_x1 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2_x1.ext -        technology: scmos
m00 w1  b z   vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=0.695475p ps=5.15u 
m01 vdd a w1  vdd p w=2.145u l=0.13u ad=1.04033p  pd=5.26u  as=0.332475p ps=2.455u
m02 z   b vss vss n w=0.605u l=0.13u ad=0.160325p pd=1.135u as=0.293425p ps=2.18u 
m03 vss a z   vss n w=0.605u l=0.13u ad=0.293425p pd=2.18u  as=0.160325p ps=1.135u
C0  a  z   0.012f
C1  a  w1  0.010f
C2  b  vdd 0.010f
C3  a  vdd 0.066f
C4  z  vdd 0.009f
C5  w1 vdd 0.010f
C6  b  a   0.196f
C7  b  z   0.081f
C9  w1 vss 0.014f
C10 z  vss 0.150f
C11 a  vss 0.125f
C12 b  vss 0.143f
.ends
