* Spice description of vfeed5
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:36
* vxlib 0.13um values
.subckt vfeed5 vdd vss
.ends
