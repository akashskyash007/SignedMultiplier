.subckt oai22v0x2 a1 a2 b1 b2 vdd vss z
*01-JAN-08 SPICE3       file   created      from oai22v0x2.ext -        technology: scmos
m00 w1  b1 vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u    as=0.635731p ps=3.17u    
m01 z   b2 w1  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u     as=0.19635p  ps=1.795u   
m02 w2  b2 z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u    as=0.3234p   ps=1.96u    
m03 vdd b1 w2  vdd p w=1.54u  l=0.13u ad=0.635731p pd=3.17u     as=0.19635p  ps=1.795u   
m04 w3  a1 vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u    as=0.635731p ps=3.17u    
m05 z   a2 w3  vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u     as=0.19635p  ps=1.795u   
m06 w4  a2 z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u    as=0.3234p   ps=1.96u    
m07 vdd a1 w4  vdd p w=1.54u  l=0.13u ad=0.635731p pd=3.17u     as=0.19635p  ps=1.795u   
m08 z   b1 n3  vss n w=0.77u  l=0.13u ad=0.1617p   pd=1.19u     as=0.18329p  ps=1.53314u 
m09 n3  b2 z   vss n w=0.77u  l=0.13u ad=0.18329p  pd=1.53314u  as=0.1617p   ps=1.19u    
m10 z   b2 n3  vss n w=0.77u  l=0.13u ad=0.1617p   pd=1.19u     as=0.18329p  ps=1.53314u 
m11 n3  b1 z   vss n w=0.77u  l=0.13u ad=0.18329p  pd=1.53314u  as=0.1617p   ps=1.19u    
m12 vss a1 n3  vss n w=0.77u  l=0.13u ad=0.255607p pd=1.81696u  as=0.18329p  ps=1.53314u 
m13 n3  a2 vss vss n w=0.77u  l=0.13u ad=0.18329p  pd=1.53314u  as=0.255607p ps=1.81696u 
m14 vss a2 n3  vss n w=0.495u l=0.13u ad=0.164318p pd=1.16804u  as=0.117829p ps=0.985588u
m15 n3  a1 vss vss n w=0.495u l=0.13u ad=0.117829p pd=0.985588u as=0.164318p ps=1.16804u 
C0  b1  w2  0.006f
C1  b2  z   0.075f
C2  vdd w4  0.004f
C3  a1  z   0.098f
C4  a2  z   0.015f
C5  vdd b1  0.022f
C6  b1  n3  0.022f
C7  a1  w3  0.006f
C8  w1  z   0.009f
C9  vdd b2  0.014f
C10 b2  n3  0.012f
C11 a1  w4  0.014f
C12 vdd a1  0.061f
C13 a1  n3  0.029f
C14 z   w2  0.009f
C15 vdd a2  0.014f
C16 b1  b2  0.333f
C17 a2  n3  0.049f
C18 z   w3  0.009f
C19 vdd w1  0.004f
C20 b1  a1  0.070f
C21 vdd z   0.132f
C22 z   n3  0.191f
C23 b1  w1  0.006f
C24 vdd w2  0.004f
C25 b1  z   0.220f
C26 vdd w3  0.004f
C27 a1  a2  0.308f
C28 n3  vss 0.417f
C29 w4  vss 0.007f
C30 w3  vss 0.007f
C31 w2  vss 0.009f
C32 z   vss 0.211f
C33 w1  vss 0.008f
C34 a2  vss 0.152f
C35 a1  vss 0.176f
C36 b2  vss 0.125f
C37 b1  vss 0.171f
.ends
