.subckt bf1_x8 a vdd vss z
*04-JAN-08 SPICE3       file   created      from bf1_x8.ext -        technology: scmos
m00 z   an vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.87793u as=0.715753p ps=3.65182u
m01 vdd an z   vdd p w=2.145u l=0.13u ad=0.715753p pd=3.65182u as=0.568425p ps=2.87793u
m02 z   an vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.87793u as=0.715753p ps=3.65182u
m03 vdd an z   vdd p w=1.54u  l=0.13u ad=0.513874p pd=2.62182u as=0.4081p   ps=2.06621u
m04 an  a  vdd vdd p w=1.54u  l=0.13u ad=0.4081p   pd=2.19625u as=0.513874p ps=2.62182u
m05 vdd a  an  vdd p w=1.98u  l=0.13u ad=0.660695p pd=3.37091u as=0.5247p   ps=2.82375u
m06 z   an vss vss n w=0.99u  l=0.13u ad=0.26235p  pd=1.52u    as=0.327271p ps=2.01635u
m07 vss an z   vss n w=0.99u  l=0.13u ad=0.327271p pd=2.01635u as=0.26235p  ps=1.52u   
m08 z   an vss vss n w=0.99u  l=0.13u ad=0.26235p  pd=1.52u    as=0.327271p ps=2.01635u
m09 vss an z   vss n w=0.99u  l=0.13u ad=0.327271p pd=2.01635u as=0.26235p  ps=1.52u   
m10 an  a  vss vss n w=0.88u  l=0.13u ad=0.2332p   pd=1.41u    as=0.290908p ps=1.79231u
m11 vss a  an  vss n w=0.88u  l=0.13u ad=0.290908p pd=1.79231u as=0.2332p   ps=1.41u   
C0 vdd an  0.061f
C1 vdd z   0.110f
C2 vdd a   0.031f
C3 an  z   0.140f
C4 an  a   0.164f
C5 a   vss 0.241f
C6 z   vss 0.403f
C7 an  vss 0.492f
.ends
