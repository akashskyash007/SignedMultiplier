* Spice description of ao22_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:01:48
* sxlib 0.13um values
.subckt ao22_x2 i0 i1 i2 q vdd vss
Mtr_00001 sig2  i0    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 sig3  i1    sig2  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 vss   i2    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00004 q     sig2  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00005 vdd   sig2  q     vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
Mtr_00006 sig2  i2    vdd   vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00007 vdd   i0    sig9  vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00008 sig9  i1    sig2  vdd p  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
C6  i0    vss   0.828f
C7  i1    vss   0.908f
C8  i2    vss   1.051f
C4  q     vss   0.944f
C2  sig2  vss   0.883f
C3  sig3  vss   0.182f
.ends
