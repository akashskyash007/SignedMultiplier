* Spice description of vfeed5
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:52
* vsclib 0.13um values
.subckt vfeed5 vdd vss
.ends
