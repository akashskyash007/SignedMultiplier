.subckt nao2o22_x1 i0 i1 i2 i3 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nao2o22_x1.ext -        technology: scmos
m00 w1  i0 vdd vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.8763p  ps=5.23u 
m01 nq  i1 w1  vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.58035p ps=2.72u 
m02 w2  i3 nq  vdd p w=2.19u l=0.13u ad=0.58035p pd=2.72u  as=0.58035p ps=2.72u 
m03 vdd i2 w2  vdd p w=2.19u l=0.13u ad=0.8763p  pd=5.23u  as=0.58035p ps=2.72u 
m04 nq  i0 w3  vss n w=1.09u l=0.13u ad=0.35925p pd=2.06u  as=0.37605p ps=2.325u
m05 w3  i1 nq  vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.35925p ps=2.06u 
m06 vss i3 w3  vss n w=1.09u l=0.13u ad=0.28885p pd=1.62u  as=0.37605p ps=2.325u
m07 w3  i2 vss vss n w=1.09u l=0.13u ad=0.37605p pd=2.325u as=0.28885p ps=1.62u 
C0  i1  w1  0.052f
C1  i3  i2  0.247f
C2  i1  nq  0.132f
C3  i3  nq  0.140f
C4  i3  w2  0.052f
C5  vdd i0  0.052f
C6  i0  w3  0.005f
C7  vdd i1  0.021f
C8  i1  w3  0.005f
C9  vdd i3  0.021f
C10 i3  w3  0.014f
C11 vdd i2  0.092f
C12 i0  i1  0.221f
C13 i2  w3  0.014f
C14 vdd w1  0.019f
C15 vdd nq  0.029f
C16 i1  i3  0.096f
C17 nq  w3  0.051f
C18 vdd w2  0.019f
C19 w3  vss 0.242f
C20 w2  vss 0.015f
C21 nq  vss 0.122f
C22 w1  vss 0.015f
C23 i2  vss 0.142f
C24 i3  vss 0.146f
C25 i1  vss 0.133f
C26 i0  vss 0.132f
.ends
