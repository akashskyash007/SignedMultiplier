.subckt oan21_x2 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from oan21_x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=2.09u  l=0.13u ad=0.755013p pd=4.06917u as=0.6809p   ps=5.04u   
m01 zn  b  vdd vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.8069u  as=0.397375p ps=2.14167u
m02 w1  a2 zn  vdd p w=2.09u  l=0.13u ad=0.32395p  pd=2.4u     as=0.55385p  ps=3.4331u 
m03 vdd a1 w1  vdd p w=2.09u  l=0.13u ad=0.755013p pd=4.06917u as=0.32395p  ps=2.4u    
m04 z   zn vss vss n w=1.045u l=0.13u ad=0.403975p pd=2.95u    as=0.371271p ps=2.62057u
m05 n2  b  zn  vss n w=0.935u l=0.13u ad=0.290125p pd=1.88667u as=0.374825p ps=2.73u   
m06 vss a2 n2  vss n w=0.935u l=0.13u ad=0.33219p  pd=2.34472u as=0.290125p ps=1.88667u
m07 n2  a1 vss vss n w=0.935u l=0.13u ad=0.290125p pd=1.88667u as=0.33219p  ps=2.34472u
C0  a2  n2  0.010f
C1  a1  w1  0.012f
C2  a1  n2  0.007f
C3  vdd zn  0.050f
C4  vdd a2  0.010f
C5  b   n2  0.073f
C6  vdd a1  0.065f
C7  zn  a2  0.013f
C8  vdd z   0.015f
C9  zn  a1  0.016f
C10 zn  z   0.145f
C11 vdd w1  0.009f
C12 a2  a1  0.224f
C13 zn  b   0.151f
C14 a2  b   0.141f
C15 zn  n2  0.007f
C16 a2  w1  0.017f
C17 a1  b   0.002f
C18 n2  vss 0.127f
C19 w1  vss 0.014f
C20 b   vss 0.125f
C21 z   vss 0.125f
C22 a1  vss 0.100f
C23 a2  vss 0.142f
C24 zn  vss 0.200f
.ends
