.subckt iv1v0x4 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v0x4.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u    as=0.61985p  ps=3.885u  
m01 vdd a z   vdd p w=1.54u  l=0.13u ad=0.61985p  pd=3.885u   as=0.3234p   ps=1.96u   
m02 z   a vss vss n w=0.935u l=0.13u ad=0.20737p  pd=1.64536u as=0.370828p ps=2.8475u 
m03 vss a z   vss n w=0.605u l=0.13u ad=0.239947p pd=1.8425u  as=0.13418p  ps=1.06464u
C0 vdd z   0.092f
C1 a   vdd 0.019f
C2 a   z   0.070f
C3 z   vss 0.162f
C5 a   vss 0.172f
.ends
