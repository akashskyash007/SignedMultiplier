.subckt aon21_x1 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from aon21_x1.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.1u   l=0.13u ad=0.341917p pd=2.06111u  as=0.34595p  ps=3.06u   
m01 n2  b  zn  vdd p w=1.43u  l=0.13u ad=0.3971p   pd=2.54667u  as=0.4334p   ps=3.72u   
m02 vdd a2 n2  vdd p w=1.43u  l=0.13u ad=0.444492p pd=2.67944u  as=0.3971p   ps=2.54667u
m03 n2  a1 vdd vdd p w=1.43u  l=0.13u ad=0.3971p   pd=2.54667u  as=0.444492p ps=2.67944u
m04 vss zn z   vss n w=0.55u  l=0.13u ad=0.267793p pd=1.76207u  as=0.2002p   ps=1.96u   
m05 zn  b  vss vss n w=0.385u l=0.13u ad=0.102025p pd=0.876842u as=0.187455p ps=1.23345u
m06 w1  a2 zn  vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u     as=0.1749p   ps=1.50316u
m07 vss a1 w1  vss n w=0.66u  l=0.13u ad=0.321352p pd=2.11448u  as=0.1023p   ps=0.97u   
C0  zn  a1  0.034f
C1  vdd b   0.022f
C2  n2  a1  0.007f
C3  vdd a2  0.012f
C4  vdd zn  0.006f
C5  a1  w1  0.014f
C6  vdd z   0.029f
C7  b   a2  0.157f
C8  vdd n2  0.106f
C9  b   zn  0.085f
C10 vdd a1  0.007f
C11 b   n2  0.070f
C12 zn  z   0.052f
C13 a2  n2  0.031f
C14 a2  a1  0.190f
C15 a1  vss 0.219f
C16 n2  vss 0.044f
C17 z   vss 0.100f
C18 zn  vss 0.179f
C19 a2  vss 0.135f
C20 b   vss 0.111f
.ends
