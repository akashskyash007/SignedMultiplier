* Spice description of an4_x1
* Spice driver version 134999461
* Date  4/01/2008 at 18:49:16
* vsxlib 0.13um values
.subckt an4_x1 a b c d vdd vss z
M1a 2z    a     vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M1b vdd   b     2z    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M1c 2z    c     vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M1d vdd   d     2z    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M1z vdd   2z    z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2a vss   a     sig5  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M2b sig5  b     n2    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M2c n2    c     sig4  vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M2d sig4  d     2z    vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
M2z z     2z    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
C3  2z    vss   1.365f
C10 a     vss   0.908f
C9  b     vss   0.886f
C8  c     vss   0.881f
C7  d     vss   0.878f
C2  z     vss   0.765f
.ends
