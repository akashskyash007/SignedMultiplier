.subckt xaon21v0x05 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from xaon21v0x05.ext -        technology: scmos
m00 z   an bn  vdd p w=0.88u  l=0.13u ad=0.1848p   pd=1.3u     as=0.265467p ps=2.42667u
m01 an  bn z   vdd p w=0.88u  l=0.13u ad=0.21651p  pd=1.7131u  as=0.1848p   ps=1.3u    
m02 vdd a2 an  vdd p w=1.155u l=0.13u ad=0.393166p pd=2.55048u as=0.28417p  ps=2.24845u
m03 vdd a1 an  vdd p w=1.155u l=0.13u ad=0.393166p pd=2.55048u as=0.28417p  ps=2.24845u
m04 bn  b  vdd vdd p w=1.1u   l=0.13u ad=0.331833p pd=3.03333u as=0.374444p ps=2.42903u
m05 w1  an vss vss n w=0.55u  l=0.13u ad=0.070125p pd=0.805u   as=0.297p    ps=1.92333u
m06 z   bn w1  vss n w=0.55u  l=0.13u ad=0.1155p   pd=0.97u    as=0.070125p ps=0.805u  
m07 an  b  z   vss n w=0.55u  l=0.13u ad=0.1155p   pd=0.97u    as=0.1155p   ps=0.97u   
m08 w2  a2 an  vss n w=0.55u  l=0.13u ad=0.070125p pd=0.805u   as=0.1155p   ps=0.97u   
m09 vss a1 w2  vss n w=0.55u  l=0.13u ad=0.297p    pd=1.92333u as=0.070125p ps=0.805u  
m10 bn  b  vss vss n w=0.55u  l=0.13u ad=0.18205p  pd=1.85u    as=0.297p    ps=1.92333u
C0  vdd a2  0.007f
C1  an  bn  0.421f
C2  an  a2  0.071f
C3  vdd a1  0.002f
C4  vdd b   0.040f
C5  an  z   0.224f
C6  bn  a2  0.130f
C7  bn  z   0.098f
C8  a2  z   0.006f
C9  an  b   0.007f
C10 bn  a1  0.041f
C11 an  w1  0.003f
C12 bn  b   0.091f
C13 a2  a1  0.140f
C14 a2  b   0.036f
C15 z   b   0.006f
C16 vdd an  0.024f
C17 a2  w2  0.013f
C18 z   w1  0.009f
C19 a1  b   0.048f
C20 vdd bn  0.195f
C21 w2  vss 0.001f
C22 w1  vss 0.004f
C23 b   vss 0.269f
C24 a1  vss 0.181f
C25 z   vss 0.289f
C26 a2  vss 0.146f
C27 bn  vss 0.215f
C28 an  vss 0.180f
.ends
