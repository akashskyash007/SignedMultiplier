.subckt xor2v1x05 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from xor2v1x05.ext -        technology: scmos
m00 an  a  vdd vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.325142p ps=2.03333u
m01 z   bn an  vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.1386p   ps=1.08u   
m02 ai  b  z   vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.1386p   ps=1.08u   
m03 vdd an ai  vdd p w=0.66u l=0.13u ad=0.325142p pd=2.03333u as=0.1386p   ps=1.08u   
m04 bn  b  vdd vdd p w=0.66u l=0.13u ad=0.2112p   pd=2.07u    as=0.325142p ps=2.03333u
m05 an  a  vss vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.1903p   ps=1.59333u
m06 z   b  an  vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.0693p   ps=0.75u   
m07 ai  bn z   vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.0693p   ps=0.75u   
m08 vss an ai  vss n w=0.33u l=0.13u ad=0.1903p   pd=1.59333u as=0.0693p   ps=0.75u   
m09 bn  b  vss vss n w=0.33u l=0.13u ad=0.12375p  pd=1.41u    as=0.1903p   ps=1.59333u
C0  b   z   0.012f
C1  bn  an  0.033f
C2  b   ai  0.021f
C3  bn  z   0.036f
C4  a   an  0.052f
C5  a   z   0.007f
C6  bn  ai  0.010f
C7  an  z   0.102f
C8  an  ai  0.113f
C9  vdd b   0.045f
C10 z   ai  0.076f
C11 vdd bn  0.104f
C12 vdd a   0.006f
C13 vdd an  0.003f
C14 b   bn  0.168f
C15 b   a   0.019f
C16 bn  a   0.028f
C17 b   an  0.090f
C18 ai  vss 0.041f
C19 z   vss 0.058f
C20 an  vss 0.366f
C21 a   vss 0.147f
C22 bn  vss 0.182f
C23 b   vss 0.253f
.ends
