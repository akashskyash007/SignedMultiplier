* Spice description of iv1v8x1
* Spice driver version 134999461
* Date  1/01/2008 at 16:47:08
* wsclib 0.13um values
.subckt iv1v8x1 a vdd vss z
M01 z     a     vdd   vdd p  L=0.12U  W=0.825U AS=0.218625P AD=0.218625P PS=2.18U   PD=2.18U
M02 vss   a     z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C3  a     vss   0.567f
C2  z     vss   0.454f
.ends
