* Spice description of one_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:36:44
* ssxlib 0.13um values
.subckt one_x0 q vdd vss
Mtr_00001 q     vss   vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
C2  q     vss   0.666f
.ends
