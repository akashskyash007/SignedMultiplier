.subckt vfeed1 vdd vss
*10-JAN-08 SPICE3       file   created      from vfeed1.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 w2  vdd vdd vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 vss vdd w3  vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m03 w4  vdd vss vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0 w4 vss 0.014f
C1 w3 vss 0.014f
C2 w2 vss 0.019f
C3 w1 vss 0.019f
.ends
