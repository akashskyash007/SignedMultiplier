* Spice description of tie_x0
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:22
* wsclib 0.13um values
.subckt tie_x0 vdd vss
.ends
