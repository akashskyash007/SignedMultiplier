.subckt an2_x05 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from an2_x05.ext -        technology: scmos
m00 vdd zn z   vdd p w=0.66u l=0.13u ad=0.3685p   pd=2.47333u as=0.22935p  ps=2.18u   
m01 zn  a  vdd vdd p w=0.66u l=0.13u ad=0.1749p   pd=1.19u    as=0.3685p   ps=2.47333u
m02 vdd b  zn  vdd p w=0.66u l=0.13u ad=0.3685p   pd=2.47333u as=0.1749p   ps=1.19u   
m03 vss zn z   vss n w=0.33u l=0.13u ad=0.223575p pd=1.34625u as=0.1419p   ps=1.52u   
m04 w1  a  vss vss n w=0.55u l=0.13u ad=0.08525p  pd=0.86u    as=0.372625p ps=2.24375u
m05 zn  b  w1  vss n w=0.55u l=0.13u ad=0.2002p   pd=1.96u    as=0.08525p  ps=0.86u   
C0  a   w2  0.012f
C1  z   w3  0.013f
C2  b   w2  0.018f
C3  z   w4  0.010f
C4  vdd b   0.016f
C5  z   w2  0.018f
C6  vdd z   0.031f
C7  zn  a   0.162f
C8  w1  w2  0.002f
C9  zn  b   0.066f
C10 w5  w2  0.166f
C11 vdd w5  0.021f
C12 zn  z   0.110f
C13 a   b   0.132f
C14 w3  w2  0.166f
C15 vdd w3  0.005f
C16 zn  w1  0.010f
C17 w4  w2  0.166f
C18 b   z   0.019f
C19 vdd w2  0.033f
C20 zn  w3  0.031f
C21 zn  w4  0.013f
C22 zn  w2  0.021f
C23 a   w4  0.025f
C24 b   w3  0.010f
C25 vdd zn  0.015f
C26 w2  vss 1.045f
C27 w4  vss 0.181f
C28 w3  vss 0.175f
C29 w5  vss 0.189f
C30 z   vss 0.030f
C31 b   vss 0.071f
C32 a   vss 0.083f
C33 zn  vss 0.124f
.ends
