.subckt mx3_x4 cmd0 cmd1 i0 i1 i2 q vdd vss
*05-JAN-08 SPICE3       file   created      from mx3_x4.ext -        technology: scmos
m00 w1  i2   w2  vdd p w=1.045u l=0.13u ad=0.276925p pd=1.61757u  as=0.335426p ps=2.06964u
m01 w3  cmd1 w1  vdd p w=0.99u  l=0.13u ad=0.3663p   pd=2.24836u  as=0.26235p  ps=1.53243u
m02 w4  cmd1 vdd vdd p w=0.77u  l=0.13u ad=0.3311p   pd=2.4u      as=0.30068p  ps=1.73423u
m03 w5  w4   w3  vdd p w=1.045u l=0.13u ad=0.161975p pd=1.355u    as=0.38665p  ps=2.37327u
m04 w2  i1   w5  vdd p w=1.045u l=0.13u ad=0.335426p pd=2.06964u  as=0.161975p ps=1.355u  
m05 vdd w6   w2  vdd p w=0.99u  l=0.13u ad=0.386588p pd=2.22972u  as=0.317772p ps=1.96071u
m06 w7  cmd0 vdd vdd p w=0.99u  l=0.13u ad=0.15345p  pd=1.3u      as=0.386588p ps=2.22972u
m07 w3  i0   w7  vdd p w=0.99u  l=0.13u ad=0.3663p   pd=2.24836u  as=0.15345p  ps=1.3u    
m08 w4  cmd1 vss vss n w=0.44u  l=0.13u ad=0.1892p   pd=1.74u     as=0.194543p ps=1.32468u
m09 vdd cmd0 w6  vdd p w=0.77u  l=0.13u ad=0.30068p  pd=1.73423u  as=0.3311p   ps=2.4u    
m10 q   w3   vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u    as=0.837607p ps=4.83106u
m11 vdd w3   q   vdd p w=2.145u l=0.13u ad=0.837607p pd=4.83106u  as=0.568425p ps=2.675u  
m12 w8  i2   w9  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.19u     as=0.24145p  ps=1.70333u
m13 w3  w4   w8  vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u  as=0.1749p   ps=1.19u   
m14 w10 cmd1 w3  vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u     as=0.2959p   ps=2.03333u
m15 w9  i1   w10 vss n w=0.66u  l=0.13u ad=0.24145p  pd=1.70333u  as=0.1023p   ps=0.97u   
m16 vss cmd0 w6  vss n w=0.33u  l=0.13u ad=0.145907p pd=0.993507u as=0.1419p   ps=1.52u   
m17 vss cmd0 w9  vss n w=0.66u  l=0.13u ad=0.291814p pd=1.98701u  as=0.24145p  ps=1.70333u
m18 w11 w6   vss vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u     as=0.291814p ps=1.98701u
m19 w3  i0   w11 vss n w=0.66u  l=0.13u ad=0.2959p   pd=2.03333u  as=0.1023p   ps=0.97u   
m20 q   w3   vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.58821u  as=0.462039p ps=3.1461u 
m21 vss w3   q   vss n w=1.1u   l=0.13u ad=0.486357p pd=3.31169u  as=0.2915p   ps=1.6718u 
C0  w4   w3   0.058f
C1  w9   w10  0.010f
C2  w2   w5   0.010f
C3  vdd  q    0.080f
C4  w6   i0   0.153f
C5  w4   i1   0.113f
C6  w4   w2   0.007f
C7  w3   q    0.149f
C8  w6   vdd  0.010f
C9  cmd0 i0   0.213f
C10 vdd  i2   0.010f
C11 w3   w9   0.057f
C12 w6   w3   0.151f
C13 cmd0 vdd  0.010f
C14 vdd  cmd1 0.049f
C15 i1   w9   0.007f
C16 i1   w6   0.091f
C17 i1   i2   0.009f
C18 i0   vdd  0.010f
C19 cmd0 w3   0.140f
C20 w3   cmd1 0.023f
C21 w2   i2   0.007f
C22 i1   cmd0 0.007f
C23 i1   cmd1 0.078f
C24 i0   w3   0.038f
C25 w2   cmd1 0.058f
C26 vdd  w3   0.102f
C27 w4   w9   0.056f
C28 i1   vdd  0.010f
C29 w4   i2   0.102f
C30 vdd  w2   0.169f
C31 i1   w3   0.060f
C32 w4   cmd1 0.232f
C33 w3   w2   0.085f
C34 vdd  w1   0.017f
C35 i1   w2   0.007f
C36 w6   w9   0.010f
C37 vdd  w5   0.010f
C38 w9   i2   0.007f
C39 w4   vdd  0.010f
C40 w9   w8   0.018f
C41 w2   w1   0.018f
C42 vdd  w7   0.010f
C43 w9   cmd1 0.007f
C44 w6   cmd0 0.252f
C45 w6   cmd1 0.005f
C46 i2   cmd1 0.114f
C47 w11  vss  0.012f
C48 w10  vss  0.008f
C49 w8   vss  0.015f
C50 w9   vss  0.218f
C51 q    vss  0.160f
C52 w7   vss  0.006f
C53 w5   vss  0.005f
C54 w1   vss  0.009f
C55 w2   vss  0.060f
C56 w3   vss  0.491f
C58 i0   vss  0.191f
C59 cmd0 vss  0.265f
C60 w6   vss  0.220f
C61 i1   vss  0.139f
C62 w4   vss  0.202f
C63 cmd1 vss  0.304f
C64 i2   vss  0.130f
.ends
