* Spice description of oa22_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:30:01
* ssxlib 0.13um values
.subckt oa22_x2 i0 i1 i2 q vdd vss
Mtr_00001 q     sig1  vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
Mtr_00002 vss   i2    sig1  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
Mtr_00003 sig3  i0    vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00004 sig1  i1    sig3  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
Mtr_00005 vdd   sig1  q     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00006 sig9  i2    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00007 sig9  i0    sig1  vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00008 sig1  i1    sig9  vdd p  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C5  i0    vss   0.807f
C4  i1    vss   0.697f
C7  i2    vss   1.025f
C6  q     vss   0.873f
C1  sig1  vss   0.835f
C9  sig9  vss   0.268f
.ends
