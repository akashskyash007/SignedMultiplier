.subckt iv1v1x8 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v1x8.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u  l=0.13u ad=0.329915p pd=2.11077u  as=0.440677p ps=2.88077u
m01 vdd a z   vdd p w=1.54u  l=0.13u ad=0.440677p pd=2.88077u  as=0.329915p ps=2.11077u
m02 z   a vdd vdd p w=1.54u  l=0.13u ad=0.329915p pd=2.11077u  as=0.440677p ps=2.88077u
m03 vdd a z   vdd p w=1.1u   l=0.13u ad=0.314769p pd=2.05769u  as=0.235654p ps=1.50769u
m04 z   a vss vss n w=0.495u l=0.13u ad=0.10829p  pd=0.793044u as=0.146168p ps=1.02261u
m05 vss a z   vss n w=1.1u   l=0.13u ad=0.324819p pd=2.27246u  as=0.240645p ps=1.76232u
m06 z   a vss vss n w=1.1u   l=0.13u ad=0.240645p pd=1.76232u  as=0.324819p ps=2.27246u
m07 vss a z   vss n w=1.1u   l=0.13u ad=0.324819p pd=2.27246u  as=0.240645p ps=1.76232u
C0 a   z   0.200f
C1 vdd a   0.050f
C2 vdd z   0.044f
C3 z   vss 0.222f
C4 a   vss 0.273f
.ends
