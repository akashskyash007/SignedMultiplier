.subckt xaon21_x05 a1 a2 b vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon21_x05.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.1u   l=0.13u ad=0.4125p   pd=2.21667u as=0.30965p  ps=2.10667u
m01 an  a2 vdd vdd p w=1.1u   l=0.13u ad=0.30965p  pd=2.10667u as=0.4125p   ps=2.21667u
m02 z   bn an  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.30965p  ps=2.10667u
m03 bn  an z   vdd p w=1.1u   l=0.13u ad=0.300575p pd=1.74u    as=0.2915p   ps=1.63u   
m04 vdd b  bn  vdd p w=1.1u   l=0.13u ad=0.4125p   pd=2.21667u as=0.300575p ps=1.74u   
m05 w1  a1 vss vss n w=0.66u  l=0.13u ad=0.1023p   pd=0.97u    as=0.52822p  ps=3.188u  
m06 an  a2 w1  vss n w=0.66u  l=0.13u ad=0.188513p pd=1.355u   as=0.1023p   ps=0.97u   
m07 z   b  an  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.36u    as=0.188513p ps=1.355u  
m08 w2  bn z   vss n w=0.495u l=0.13u ad=0.076725p pd=0.805u   as=0.131175p ps=1.02u   
m09 vss an w2  vss n w=0.495u l=0.13u ad=0.396165p pd=2.391u   as=0.076725p ps=0.805u  
m10 bn  b  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.396165p ps=2.391u  
C0  w3  z   0.022f
C1  w4  an  0.015f
C2  w5  w3  0.166f
C3  w3  w1  0.005f
C4  w6  a1  0.002f
C5  a1  an  0.014f
C6  a2  bn  0.039f
C7  w4  b   0.004f
C8  w3  w2  0.003f
C9  w6  a2  0.002f
C10 a2  an  0.064f
C11 w4  z   0.019f
C12 w6  bn  0.017f
C13 w3  vdd 0.057f
C14 a1  z   0.016f
C15 a2  b   0.023f
C16 bn  an  0.257f
C17 w6  an  0.008f
C18 w5  a1  0.010f
C19 a2  z   0.083f
C20 a1  w1  0.005f
C21 bn  b   0.137f
C22 w4  w3  0.166f
C23 w6  b   0.001f
C24 w3  a1  0.030f
C25 w5  a2  0.013f
C26 bn  z   0.020f
C27 an  b   0.136f
C28 w4  vdd 0.002f
C29 w6  z   0.004f
C30 w3  a2  0.018f
C31 w5  bn  0.011f
C32 an  z   0.214f
C33 w3  bn  0.028f
C34 w5  an  0.010f
C35 b   z   0.008f
C36 vdd a2  0.013f
C37 w6  w3  0.166f
C38 w4  a1  0.002f
C39 w3  an  0.082f
C40 w5  b   0.011f
C41 an  w2  0.006f
C42 vdd bn  0.084f
C43 w4  a2  0.030f
C44 w3  b   0.048f
C45 w5  z   0.009f
C46 w6  vdd 0.027f
C47 vdd an  0.045f
C48 a1  a2  0.098f
C49 w4  bn  0.011f
C50 w3  vss 0.954f
C51 w5  vss 0.174f
C52 w4  vss 0.166f
C53 w6  vss 0.168f
C54 z   vss 0.027f
C55 b   vss 0.329f
C56 an  vss 0.184f
C57 bn  vss 0.119f
C58 a2  vss 0.099f
C59 a1  vss 0.116f
.ends
