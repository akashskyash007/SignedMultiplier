.subckt nd2_x1 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nd2_x1.ext -        technology: scmos
m00 z   b vdd vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u  as=0.5335p   ps=3.17u 
m01 vdd a z   vdd p w=1.1u   l=0.13u ad=0.5335p   pd=3.17u  as=0.2915p   ps=1.63u 
m02 w1  b z   vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u as=0.374825p ps=2.73u 
m03 vss a w1  vss n w=0.935u l=0.13u ad=0.453475p pd=2.84u  as=0.144925p ps=1.245u
C0 vdd b   0.008f
C1 vdd z   0.064f
C2 b   a   0.160f
C3 b   z   0.081f
C4 a   z   0.016f
C5 a   w1  0.012f
C6 w1  vss 0.006f
C7 z   vss 0.112f
C8 a   vss 0.140f
C9 b   vss 0.117f
.ends
