* Spice description of rowend_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:36:56
* sxlib 0.13um values
.subckt rowend_x0 vdd vss
.ends
