.subckt xor2v8x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from xor2v8x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u l=0.13u ad=0.551031p pd=3.71875u as=0.4444p   ps=3.83u   
m01 bn  b  vdd vdd p w=0.66u l=0.13u ad=0.2112p   pd=2.07u    as=0.236156p ps=1.59375u
m02 an  a  vdd vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.236156p ps=1.59375u
m03 zn  b  an  vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.1386p   ps=1.08u   
m04 ai  bn zn  vdd p w=0.66u l=0.13u ad=0.1386p   pd=1.08u    as=0.1386p   ps=1.08u   
m05 vdd an ai  vdd p w=0.66u l=0.13u ad=0.236156p pd=1.59375u as=0.1386p   ps=1.08u   
m06 vss zn z   vss n w=0.77u l=0.13u ad=0.384038p pd=2.99688u as=0.24035p  ps=2.29u   
m07 an  a  vss vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.164588p ps=1.28438u
m08 zn  bn an  vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.0693p   ps=0.75u   
m09 ai  b  zn  vss n w=0.33u l=0.13u ad=0.0693p   pd=0.75u    as=0.0693p   ps=0.75u   
m10 vss an ai  vss n w=0.33u l=0.13u ad=0.164588p pd=1.28438u as=0.0693p   ps=0.75u   
m11 bn  b  vss vss n w=0.33u l=0.13u ad=0.12375p  pd=1.41u    as=0.164588p ps=1.28438u
C0  bn  an  0.140f
C1  vdd z   0.012f
C2  bn  ai  0.008f
C3  vdd b   0.039f
C4  an  ai  0.090f
C5  zn  z   0.062f
C6  vdd a   0.072f
C7  zn  b   0.006f
C8  vdd bn  0.102f
C9  vdd an  0.023f
C10 zn  a   0.066f
C11 z   a   0.023f
C12 zn  bn  0.015f
C13 zn  an  0.163f
C14 b   a   0.037f
C15 zn  ai  0.081f
C16 z   an  0.007f
C17 b   bn  0.143f
C18 a   bn  0.025f
C19 b   an  0.095f
C20 a   an  0.010f
C21 b   ai  0.020f
C22 vdd zn  0.007f
C23 ai  vss 0.029f
C24 an  vss 0.150f
C25 bn  vss 0.137f
C26 a   vss 0.087f
C27 b   vss 0.357f
C28 z   vss 0.097f
C29 zn  vss 0.254f
.ends
