.subckt iv1v5x8 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v5x8.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u l=0.13u ad=0.329915p pd=2.11077u as=0.440677p ps=2.88077u
m01 vdd a z   vdd p w=1.54u l=0.13u ad=0.440677p pd=2.88077u as=0.329915p ps=2.11077u
m02 z   a vdd vdd p w=1.54u l=0.13u ad=0.329915p pd=2.11077u as=0.440677p ps=2.88077u
m03 vdd a z   vdd p w=1.1u  l=0.13u ad=0.314769p pd=2.05769u as=0.235654p ps=1.50769u
m04 z   a vss vss n w=1.1u  l=0.13u ad=0.231p    pd=1.52u    as=0.473p    ps=3.06u   
m05 vss a z   vss n w=1.1u  l=0.13u ad=0.473p    pd=3.06u    as=0.231p    ps=1.52u   
C0 vdd a   0.021f
C1 vdd z   0.071f
C2 a   z   0.128f
C3 z   vss 0.155f
C4 a   vss 0.248f
.ends
