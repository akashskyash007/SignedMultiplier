.subckt oa2a2a2a24_x4 i0 i1 i2 i3 i4 i5 i6 i7 q vdd vss
*05-JAN-08 SPICE3       file   created      from oa2a2a2a24_x4.ext -        technology: scmos
m00 w1  i7 w2  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.726275p ps=3.83u   
m01 w2  i6 w1  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.55385p  ps=2.62u   
m02 w2  i5 w3  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.726275p ps=3.83u   
m03 w3  i4 w2  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.726275p ps=3.83u   
m04 w4  i3 w3  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.726275p ps=3.83u   
m05 w3  i2 w4  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83u    as=0.55385p  ps=2.62u   
m06 w4  i1 vdd vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.726275p ps=3.83455u
m07 vdd i0 w4  vdd p w=2.09u  l=0.13u ad=0.726275p pd=3.83455u as=0.55385p  ps=2.62u   
m08 q   w1 vdd vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.745388p ps=3.93545u
m09 vdd w1 q   vdd p w=2.145u l=0.13u ad=0.745388p pd=3.93545u as=0.568425p ps=2.675u  
m10 w5  i7 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.392892p ps=2.51372u
m11 w1  i6 w5  vss n w=1.045u l=0.13u ad=0.361988p pd=2.2648u  as=0.276925p ps=1.575u  
m12 w6  i5 vss vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.392892p ps=2.51372u
m13 w1  i4 w6  vss n w=1.045u l=0.13u ad=0.361988p pd=2.2648u  as=0.161975p ps=1.355u  
m14 w7  i3 w1  vss n w=1.045u l=0.13u ad=0.161975p pd=1.355u   as=0.361988p ps=2.2648u 
m15 vss i2 w7  vss n w=1.045u l=0.13u ad=0.392892p pd=2.51372u as=0.161975p ps=1.355u  
m16 w8  i1 w1  vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.342936p ps=2.1456u 
m17 vss i0 w8  vss n w=0.99u  l=0.13u ad=0.372214p pd=2.38142u as=0.15345p  ps=1.3u    
m18 q   w1 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u   as=0.392892p ps=2.51372u
m19 vss w1 q   vss n w=1.045u l=0.13u ad=0.392892p pd=2.51372u as=0.276925p ps=1.575u  
C0  i5  i4  0.232f
C1  w2  w3  0.097f
C2  i0  vdd 0.060f
C3  i5  w1  0.019f
C4  i3  i2  0.232f
C5  i7  i6  0.096f
C6  i4  vdd 0.010f
C7  i0  q   0.119f
C8  w1  vdd 0.037f
C9  i5  w2  0.028f
C10 w1  q   0.007f
C11 w3  w4  0.088f
C12 w2  vdd 0.122f
C13 i5  w3  0.007f
C14 i4  i3  0.200f
C15 w1  w5  0.015f
C16 w3  vdd 0.190f
C17 i3  w1  0.019f
C18 w1  i7  0.117f
C19 i5  vdd 0.010f
C20 w1  w6  0.010f
C21 w4  vdd 0.097f
C22 i2  w1  0.024f
C23 i1  i0  0.121f
C24 w1  i6  0.112f
C25 w2  i7  0.016f
C26 w1  w7  0.010f
C27 i3  w3  0.016f
C28 i1  w1  0.069f
C29 w2  i6  0.037f
C30 vdd q   0.083f
C31 i2  w3  0.007f
C32 i0  w1  0.119f
C33 i4  w1  0.019f
C34 i2  w4  0.034f
C35 i3  vdd 0.010f
C36 vdd i7  0.010f
C37 i4  w2  0.005f
C38 i1  w4  0.019f
C39 w1  w2  0.059f
C40 i2  vdd 0.010f
C41 vdd i6  0.010f
C42 i4  w3  0.012f
C43 i0  w4  0.010f
C44 i1  vdd 0.019f
C45 w8  vss 0.017f
C46 w7  vss 0.014f
C47 w6  vss 0.014f
C48 w5  vss 0.025f
C49 q   vss 0.149f
C51 w4  vss 0.068f
C52 w3  vss 0.107f
C53 w2  vss 0.125f
C54 w1  vss 0.814f
C55 i0  vss 0.137f
C56 i1  vss 0.131f
C57 i2  vss 0.129f
C58 i3  vss 0.136f
C59 i4  vss 0.124f
C60 i5  vss 0.135f
C61 i6  vss 0.150f
C62 i7  vss 0.169f
.ends
