* Spice description of an2v2x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:34:37
* wsclib 0.13um values
.subckt an2v2x2 a b vdd vss z
M01 06    a     vdd   vdd p  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M02 n1    a     vss   vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M03 vdd   b     06    vdd p  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M04 06    b     n1    vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
M05 vdd   06    z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M06 vss   06    z     vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C4  06    vss   0.638f
C5  a     vss   0.579f
C6  b     vss   0.472f
C3  z     vss   0.708f
.ends
