.subckt oan22_x2 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from oan22_x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=2.145u l=0.13u ad=0.725725p pd=3.53667u as=0.695475p ps=5.15u   
m01 w1  b1 vdd vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u   as=0.725725p ps=3.53667u
m02 zn  b2 w1  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u   as=0.332475p ps=2.455u  
m03 w2  a2 zn  vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u   as=0.568425p ps=2.675u  
m04 vdd a1 w2  vdd p w=2.145u l=0.13u ad=0.725725p pd=3.53667u as=0.332475p ps=2.455u  
m05 z   zn vss vss n w=1.045u l=0.13u ad=0.331375p pd=2.95u    as=0.391875p ps=2.66u   
m06 zn  b1 n3  vss n w=0.935u l=0.13u ad=0.247775p pd=1.465u   as=0.29315p  ps=2.0975u 
m07 n3  b2 zn  vss n w=0.935u l=0.13u ad=0.29315p  pd=2.0975u  as=0.247775p ps=1.465u  
m08 vss a2 n3  vss n w=0.935u l=0.13u ad=0.350625p pd=2.38u    as=0.29315p  ps=2.0975u 
m09 n3  a1 vss vss n w=0.935u l=0.13u ad=0.29315p  pd=2.0975u  as=0.350625p ps=2.38u   
C0  a1  n3  0.007f
C1  zn  b2  0.019f
C2  vdd a1  0.052f
C3  vdd z   0.033f
C4  b1  b2  0.197f
C5  b1  a2  0.019f
C6  zn  a1  0.019f
C7  vdd w1  0.010f
C8  zn  z   0.136f
C9  vdd w2  0.010f
C10 b2  a2  0.166f
C11 zn  w1  0.010f
C12 b2  a1  0.003f
C13 b1  w1  0.014f
C14 a2  a1  0.230f
C15 zn  n3  0.066f
C16 vdd zn  0.093f
C17 b1  n3  0.007f
C18 vdd b1  0.010f
C19 a2  w2  0.010f
C20 b2  n3  0.081f
C21 vdd b2  0.010f
C22 a2  n3  0.010f
C23 a1  w2  0.013f
C24 vdd a2  0.010f
C25 zn  b1  0.225f
C26 n3  vss 0.227f
C27 w2  vss 0.009f
C28 w1  vss 0.009f
C29 z   vss 0.116f
C30 a1  vss 0.101f
C31 a2  vss 0.116f
C32 b2  vss 0.118f
C33 b1  vss 0.123f
C34 zn  vss 0.185f
.ends
