* Spice description of aoi21v0x1
* Spice driver version 134999461
* Date  1/01/2008 at 16:37:23
* vsclib 0.13um values
.subckt aoi21v0x1 a1 a2 b vdd vss z
M01 03    a1    vdd   vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M02 vss   a1    sig3  vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M03 vdd   a2    03    vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M04 sig3  a2    z     vss n  L=0.12U  W=0.66U  AS=0.1749P   AD=0.1749P   PS=1.85U   PD=1.85U
M05 03    b     z     vdd p  L=0.12U  W=1.485U AS=0.393525P AD=0.393525P PS=3.5U    PD=3.5U
M06 z     b     vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C8  03    vss   0.291f
C4  a1    vss   0.482f
C5  a2    vss   0.459f
C6  b     vss   0.588f
C2  z     vss   0.794f
.ends
