.subckt xnr2v0x1 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from xnr2v0x1.ext -        technology: scmos
m00 vdd vdd w1  vdd p w=1.54u l=0.13u ad=0.54725p pd=3.28u as=0.5775p  ps=3.83u
m01 w2  b   vdd vdd p w=1.54u l=0.13u ad=0.5775p  pd=3.83u as=0.54725p ps=3.28u
m02 w3  w4  vdd vdd p w=1.54u l=0.13u ad=0.517p   pd=2.73u as=0.54725p ps=3.28u
m03 z   w2  w3  vdd p w=1.54u l=0.13u ad=0.5775p  pd=3.83u as=0.517p   ps=2.73u
m04 w4  b   z   vdd p w=1.54u l=0.13u ad=0.517p   pd=2.73u as=0.5775p  ps=3.83u
m05 vdd a   w4  vdd p w=1.54u l=0.13u ad=0.54725p pd=3.28u as=0.517p   ps=2.73u
m06 vss vdd w5  vss n w=1.1u  l=0.13u ad=0.4004p  pd=2.29u as=0.4125p  ps=2.95u
m07 w2  b   vss vss n w=1.1u  l=0.13u ad=0.4125p  pd=2.95u as=0.4004p  ps=2.29u
m08 z   w4  w2  vss n w=1.1u  l=0.13u ad=0.4004p  pd=2.29u as=0.4125p  ps=2.95u
m09 w4  w2  z   vss n w=1.1u  l=0.13u ad=0.4125p  pd=2.95u as=0.4004p  ps=2.29u
m10 vss b   w2  vss n w=1.1u  l=0.13u ad=0.4004p  pd=2.29u as=0.4125p  ps=2.95u
m11 w4  a   vss vss n w=1.1u  l=0.13u ad=0.4125p  pd=2.95u as=0.4004p  ps=2.29u
C0  w4  z   0.256f
C1  w3  z   0.020f
C2  vdd b   0.384f
C3  w2  z   0.067f
C4  vdd w4  0.037f
C5  vdd w3  0.008f
C6  vdd w2  0.023f
C7  b   w4  0.090f
C8  b   w3  0.010f
C9  vdd a   0.038f
C10 w4  w3  0.017f
C11 b   w2  0.106f
C12 b   a   0.089f
C13 w4  w2  0.240f
C14 w4  a   0.108f
C15 b   z   0.028f
C16 w5  vss 0.014f
C17 z   vss 0.116f
C18 w1  vss 0.019f
C19 a   vss 0.155f
C20 w2  vss 0.306f
C21 w3  vss 0.019f
C22 w4  vss 0.307f
C23 b   vss 0.322f
.ends
