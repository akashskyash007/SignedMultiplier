.subckt xnr2_x05 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from xnr2_x05.ext -        technology: scmos
m00 w1  an vdd vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u    as=0.420567p ps=2.43667u
m01 z   bn w1  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.1705p   ps=1.41u   
m02 an  b  z   vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.2915p   ps=1.63u   
m03 vdd a  an  vdd p w=1.1u   l=0.13u ad=0.420567p pd=2.43667u as=0.2915p   ps=1.63u   
m04 bn  b  vdd vdd p w=1.1u   l=0.13u ad=0.41855p  pd=3.06u    as=0.420567p ps=2.43667u
m05 z   an bn  vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u   as=0.185625p ps=1.85u   
m06 an  bn z   vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u   as=0.131175p ps=1.025u  
m07 vss a  an  vss n w=0.495u l=0.13u ad=0.6787p   pd=2.51u    as=0.131175p ps=1.025u  
m08 bn  b  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.6787p   ps=2.51u   
C0  b   w2  0.015f
C1  a   w3  0.015f
C2  z   w4  0.028f
C3  vdd a   0.004f
C4  an  bn  0.226f
C5  a   w2  0.033f
C6  z   w5  0.009f
C7  an  b   0.084f
C8  z   w3  0.030f
C9  vdd z   0.082f
C10 bn  b   0.173f
C11 z   w2  0.030f
C12 vdd w4  0.017f
C13 bn  a   0.182f
C14 w4  w2  0.166f
C15 an  z   0.169f
C16 b   a   0.134f
C17 w5  w2  0.166f
C18 an  w4  0.016f
C19 bn  z   0.044f
C20 w3  w2  0.166f
C21 vdd w2  0.050f
C22 an  w5  0.011f
C23 bn  w4  0.007f
C24 b   z   0.004f
C25 an  w3  0.009f
C26 bn  w5  0.013f
C27 b   w4  0.013f
C28 vdd an  0.015f
C29 an  w2  0.038f
C30 bn  w3  0.021f
C31 b   w5  0.043f
C32 a   w4  0.002f
C33 w1  z   0.024f
C34 vdd bn  0.010f
C35 bn  w2  0.071f
C36 b   w3  0.002f
C37 w1  w4  0.002f
C38 vdd b   0.056f
C39 w2  vss 0.981f
C40 w3  vss 0.171f
C41 w5  vss 0.170f
C42 w4  vss 0.159f
C43 z   vss 0.040f
C44 a   vss 0.180f
C45 b   vss 0.123f
C46 bn  vss 0.296f
C47 an  vss 0.112f
.ends
