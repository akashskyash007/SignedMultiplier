.subckt cgi2a_x05 a b c vdd vss z
*04-JAN-08 SPICE3       file   created      from cgi2a_x05.ext -        technology: scmos
m00 vdd b  n2  vdd p w=1.1u   l=0.13u ad=0.304163p pd=1.66977u as=0.33385p  ps=2.10667u
m01 w1  b  vdd vdd p w=1.1u   l=0.13u ad=0.1705p   pd=1.41u    as=0.304163p ps=1.66977u
m02 z   an w1  vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.1705p   ps=1.41u   
m03 n2  c  z   vdd p w=1.1u   l=0.13u ad=0.33385p  pd=2.10667u as=0.2915p   ps=1.63u   
m04 vdd an n2  vdd p w=1.1u   l=0.13u ad=0.304163p pd=1.66977u as=0.33385p  ps=2.10667u
m05 an  a  vdd vdd p w=1.43u  l=0.13u ad=0.4334p   pd=3.72u    as=0.395412p ps=2.1707u 
m06 vss b  n4  vss n w=0.495u l=0.13u ad=0.23463p  pd=1.764u   as=0.149325p ps=1.3u    
m07 w2  b  vss vss n w=0.495u l=0.13u ad=0.076725p pd=0.805u   as=0.23463p  ps=1.764u  
m08 z   an w2  vss n w=0.495u l=0.13u ad=0.131175p pd=1.025u   as=0.076725p ps=0.805u  
m09 n4  c  z   vss n w=0.495u l=0.13u ad=0.149325p pd=1.3u     as=0.131175p ps=1.025u  
m10 vss an n4  vss n w=0.495u l=0.13u ad=0.23463p  pd=1.764u   as=0.149325p ps=1.3u    
m11 an  a  vss vss n w=0.715u l=0.13u ad=0.243925p pd=2.29u    as=0.33891p  ps=2.548u  
C0  w3  w4  0.166f
C1  w4  w1  0.002f
C2  w5  z   0.009f
C3  w2  w4  0.002f
C4  w3  vdd 0.026f
C5  an  c   0.211f
C6  w6  w4  0.166f
C7  w4  z   0.023f
C8  w6  vdd 0.004f
C9  b   n2  0.027f
C10 an  a   0.166f
C11 n4  z   0.052f
C12 w5  w4  0.166f
C13 w3  b   0.005f
C14 c   a   0.067f
C15 an  n2  0.007f
C16 w4  vdd 0.049f
C17 w6  b   0.012f
C18 w3  an  0.008f
C19 b   z   0.016f
C20 c   n2  0.040f
C21 n4  w4  0.061f
C22 w3  c   0.001f
C23 w5  b   0.013f
C24 w6  an  0.014f
C25 an  z   0.092f
C26 w4  b   0.023f
C27 w5  an  0.071f
C28 w6  c   0.011f
C29 w3  a   0.002f
C30 c   z   0.073f
C31 vdd b   0.004f
C32 n4  b   0.011f
C33 w4  an  0.032f
C34 w6  a   0.011f
C35 w3  n2  0.043f
C36 n2  w1  0.029f
C37 vdd an  0.004f
C38 n4  an  0.018f
C39 w4  c   0.016f
C40 w3  w1  0.002f
C41 n2  z   0.056f
C42 vdd c   0.002f
C43 n4  c   0.005f
C44 w3  z   0.005f
C45 w4  a   0.026f
C46 w1  z   0.001f
C47 w2  z   0.012f
C48 vdd a   0.053f
C49 b   an  0.135f
C50 w4  n2  0.023f
C51 w6  z   0.030f
C52 vdd n2  0.146f
C53 w4  vss 0.967f
C54 w5  vss 0.165f
C55 w6  vss 0.167f
C56 w3  vss 0.154f
C57 n4  vss 0.175f
C58 z   vss 0.030f
C59 n2  vss 0.002f
C60 a   vss 0.069f
C61 c   vss 0.091f
C62 an  vss 0.191f
C63 b   vss 0.172f
.ends
