* Spice description of vfeed3
* Spice driver version 134999461
* Date  4/01/2008 at 19:51:25
* vsxlib 0.13um values
.subckt vfeed3 vdd vss
.ends
