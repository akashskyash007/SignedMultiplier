* Spice description of nr2av0x1
* Spice driver version 134999461
* Date 10/01/2008 at 14:51:09
* rgalib 0.13um values
.subckt nr2av0x1 a b vdd vss z
Mtr_00001 vss   vdd   sig3  vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00002 sig1  a     vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00003 z     sig1  vss   vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00004 vss   b     z     vss n  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00005 vdd   vdd   sig8  vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00006 sig1  a     vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00007 sig9  sig1  vdd   vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
Mtr_00008 z     b     sig9  vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
C5  a     vss   0.602f
C7  b     vss   0.558f
C1  sig1  vss   0.755f
C6  z     vss   0.644f
.ends
