.subckt na2_x4 i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from na2_x4.ext -        technology: scmos
m00 w1  i0 vdd vdd p w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.358054p ps=2.10733u
m01 vdd i1 w1  vdd p w=1.09u l=0.13u ad=0.358054p pd=2.10733u as=0.28885p  ps=1.62u   
m02 nq  w2 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.719394p ps=4.234u  
m03 vdd w2 nq  vdd p w=2.19u l=0.13u ad=0.719394p pd=4.234u   as=0.58035p  ps=2.72u   
m04 w2  w1 vdd vdd p w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.358054p ps=2.10733u
m05 w3  i0 w1  vss n w=1.09u l=0.13u ad=0.2289p   pd=1.51u    as=0.46325p  ps=3.03u   
m06 vss i1 w3  vss n w=1.09u l=0.13u ad=0.364378p pd=2.16856u as=0.2289p   ps=1.51u   
m07 nq  w2 vss vss n w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.364378p ps=2.16856u
m08 vss w2 nq  vss n w=1.09u l=0.13u ad=0.364378p pd=2.16856u as=0.28885p  ps=1.62u   
m09 w2  w1 vss vss n w=0.54u l=0.13u ad=0.2295p   pd=1.93u    as=0.180517p ps=1.07433u
C0  i1  w1  0.141f
C1  i1  w3  0.009f
C2  w1  nq  0.145f
C3  w1  w3  0.011f
C4  w2  vdd 0.020f
C5  w2  i1  0.051f
C6  vdd i0  0.011f
C7  w2  w1  0.094f
C8  vdd i1  0.002f
C9  w2  nq  0.030f
C10 vdd w1  0.168f
C11 i0  i1  0.207f
C12 i0  w1  0.023f
C13 vdd nq  0.019f
C14 w3  vss 0.008f
C15 nq  vss 0.112f
C16 w1  vss 0.280f
C17 i1  vss 0.133f
C18 i0  vss 0.128f
C20 w2  vss 0.279f
.ends
