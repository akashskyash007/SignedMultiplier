.subckt inv_x4 i nq vdd vss
*05-JAN-08 SPICE3       file   created      from inv_x4.ext -        technology: scmos
m00 nq  i vdd vdd p w=2.145u l=0.13u ad=0.632775p pd=3.16136u as=0.92235p  ps=5.30636u
m01 vdd i nq  vdd p w=1.485u l=0.13u ad=0.63855p  pd=3.67364u as=0.438075p ps=2.18864u
m02 nq  i vss vss n w=0.99u  l=0.13u ad=0.26235p  pd=1.52u    as=0.4257p   ps=2.84u   
m03 vss i nq  vss n w=0.99u  l=0.13u ad=0.4257p   pd=2.84u    as=0.26235p  ps=1.52u   
C0 vdd nq  0.061f
C1 i   vdd 0.087f
C2 i   nq  0.191f
C3 nq  vss 0.131f
C5 i   vss 0.314f
.ends
