* Spice description of vfeed3
* Spice driver version 134999461
* Date  1/01/2008 at 17:02:42
* vsclib 0.13um values
.subckt vfeed3 vdd vss
.ends
