.subckt bf1_x1 a vdd vss z
*04-JAN-08 SPICE3       file   created      from bf1_x1.ext -        technology: scmos
m00 vdd an z   vdd p w=1.1u  l=0.13u ad=0.2915p  pd=1.63u as=0.41855p ps=3.06u
m01 an  a  vdd vdd p w=1.1u  l=0.13u ad=0.41855p pd=3.06u as=0.2915p  ps=1.63u
m02 vss an z   vss n w=0.55u l=0.13u ad=0.2002p  pd=1.41u as=0.2002p  ps=1.96u
m03 an  a  vss vss n w=0.55u l=0.13u ad=0.2002p  pd=1.96u as=0.2002p  ps=1.41u
C0 vdd an  0.064f
C1 vdd a   0.002f
C2 vdd z   0.006f
C3 an  a   0.187f
C4 an  z   0.114f
C5 z   vss 0.075f
C6 a   vss 0.121f
C7 an  vss 0.197f
.ends
