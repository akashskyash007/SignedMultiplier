* Spice description of zero_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:43:45
* sxlib 0.13um values
.subckt zero_x0 nq vdd vss
Mtr_00001 vss   vdd   nq    vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
C1  nq    vss   0.704f
.ends
