.subckt an3v0x2 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from an3v0x2.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.54u  l=0.13u ad=0.422038p pd=2.66177u as=0.48675p  ps=3.83u   
m01 zn  a  vdd vdd p w=0.935u l=0.13u ad=0.225592p pd=1.77667u as=0.256237p ps=1.61608u
m02 vdd b  zn  vdd p w=0.935u l=0.13u ad=0.256237p pd=1.61608u as=0.225592p ps=1.77667u
m03 zn  c  vdd vdd p w=0.935u l=0.13u ad=0.225592p pd=1.77667u as=0.256237p ps=1.61608u
m04 vss zn z   vss n w=0.77u  l=0.13u ad=0.287384p pd=1.62129u as=0.24035p  ps=2.29u   
m05 w1  a  vss vss n w=0.935u l=0.13u ad=0.119213p pd=1.19u    as=0.348966p ps=1.96871u
m06 w2  b  w1  vss n w=0.935u l=0.13u ad=0.119213p pd=1.19u    as=0.119213p ps=1.19u   
m07 zn  c  w2  vss n w=0.935u l=0.13u ad=0.284075p pd=2.62u    as=0.119213p ps=1.19u   
C0  zn  w2  0.008f
C1  a   c   0.030f
C2  b   c   0.138f
C3  zn  z   0.152f
C4  zn  vdd 0.135f
C5  c   w2  0.005f
C6  z   vdd 0.004f
C7  zn  a   0.177f
C8  z   a   0.007f
C9  zn  b   0.034f
C10 zn  c   0.060f
C11 vdd a   0.006f
C12 vdd b   0.006f
C13 zn  w1  0.014f
C14 vdd c   0.006f
C15 a   b   0.139f
C16 w2  vss 0.007f
C17 w1  vss 0.006f
C18 c   vss 0.108f
C19 b   vss 0.100f
C20 a   vss 0.102f
C22 z   vss 0.210f
C23 zn  vss 0.245f
.ends
