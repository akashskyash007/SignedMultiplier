* Spice description of an3v4x2
* Spice driver version 134999461
* Date  1/01/2008 at 16:35:35
* vsclib 0.13um values
.subckt an3v4x2 a b c vdd vss z
M01 08    a     vdd   vdd p  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M02 n1    a     vss   vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M03 vdd   b     08    vdd p  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M04 sig7  b     n1    vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M05 08    c     vdd   vdd p  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M06 08    c     sig7  vss n  L=0.12U  W=0.495U AS=0.131175P AD=0.131175P PS=1.52U   PD=1.52U
M07 vdd   08    z     vdd p  L=0.12U  W=1.54U  AS=0.4081P   AD=0.4081P   PS=3.61U   PD=3.61U
M08 vss   08    z     vss n  L=0.12U  W=0.77U  AS=0.20405P  AD=0.20405P  PS=2.07U   PD=2.07U
C4  08    vss   0.790f
C5  a     vss   0.665f
C8  b     vss   0.687f
C6  c     vss   0.732f
C2  z     vss   0.628f
.ends
