.subckt noa22_x1 i0 i1 i2 nq vdd vss
*05-JAN-08 SPICE3       file   created      from noa22_x1.ext -        technology: scmos
m00 nq  i0 w1  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.6864p   ps=3.5u  
m01 w1  i1 nq  vdd p w=2.145u l=0.13u ad=0.6864p   pd=3.5u   as=0.568425p ps=2.675u
m02 vdd i2 w1  vdd p w=2.145u l=0.13u ad=0.92235p  pd=5.15u  as=0.6864p   ps=3.5u  
m03 w2  i0 vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u as=0.44935p  ps=2.95u 
m04 nq  i1 w2  vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u as=0.276925p ps=1.575u
m05 vss i2 nq  vss n w=1.045u l=0.13u ad=0.44935p  pd=2.95u  as=0.276925p ps=1.575u
C0  vdd i1  0.010f
C1  vdd i2  0.120f
C2  vdd w1  0.108f
C3  i0  i1  0.226f
C4  vdd nq  0.017f
C5  i1  i2  0.096f
C6  i0  w1  0.017f
C7  i1  w1  0.007f
C8  i2  w1  0.012f
C9  i1  nq  0.155f
C10 i2  nq  0.145f
C11 i1  w2  0.017f
C12 w1  nq  0.111f
C13 vdd i0  0.010f
C14 w2  vss 0.024f
C15 nq  vss 0.128f
C16 w1  vss 0.091f
C17 i2  vss 0.224f
C18 i1  vss 0.163f
C19 i0  vss 0.167f
.ends
