.subckt vfeed1 vdd vss
*01-JAN-08 SPICE3       file   created      from vfeed1.ext -        technology: scmos
.ends
