.subckt iv1v0x1 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v0x1.ext -        technology: scmos
m00 vdd a z vdd p w=0.99u  l=0.13u ad=0.543675p pd=3.28u as=0.341p    ps=2.73u
m01 vss a z vss n w=0.495u l=0.13u ad=0.294525p pd=2.18u as=0.167475p ps=1.74u
C0 vdd z   0.013f
C1 a   z   0.073f
C2 z   vss 0.184f
C3 a   vss 0.117f
.ends
