.subckt iv1_x3 a vdd vss z
*04-JAN-08 SPICE3       file   created      from iv1_x3.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u l=0.13u ad=0.4081p  pd=2.07u as=0.7469p  ps=4.05u
m01 vdd a z   vdd p w=1.54u l=0.13u ad=0.7469p  pd=4.05u as=0.4081p  ps=2.07u
m02 z   a vss vss n w=0.77u l=0.13u ad=0.20405p pd=1.3u  as=0.37345p ps=2.51u
m03 vss a z   vss n w=0.77u l=0.13u ad=0.37345p pd=2.51u as=0.20405p ps=1.3u 
C0  vdd z   0.045f
C1  vdd w1  0.025f
C2  vdd w2  0.007f
C3  a   z   0.092f
C4  a   w1  0.005f
C5  z   w1  0.008f
C6  vdd w3  0.048f
C7  a   w2  0.011f
C8  z   w2  0.033f
C9  a   w4  0.011f
C10 a   w3  0.018f
C11 z   w4  0.031f
C12 z   w3  0.020f
C13 w1  w3  0.166f
C14 w2  w3  0.166f
C15 vdd a   0.029f
C16 w4  w3  0.166f
C17 w3  vss 1.068f
C18 w4  vss 0.184f
C19 w2  vss 0.177f
C20 w1  vss 0.177f
C21 z   vss 0.069f
C22 a   vss 0.131f
.ends
