.subckt nd2v0x8 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nd2v0x8.ext -        technology: scmos
m00 z   a vdd vdd p w=1.43u l=0.13u ad=0.3003p   pd=1.885u   as=0.360926p ps=2.36167u
m01 vdd b z   vdd p w=1.43u l=0.13u ad=0.360926p pd=2.36167u as=0.3003p   ps=1.885u  
m02 z   b vdd vdd p w=1.43u l=0.13u ad=0.3003p   pd=1.885u   as=0.360926p ps=2.36167u
m03 vdd a z   vdd p w=1.43u l=0.13u ad=0.360926p pd=2.36167u as=0.3003p   ps=1.885u  
m04 z   a vdd vdd p w=1.43u l=0.13u ad=0.3003p   pd=1.885u   as=0.360926p ps=2.36167u
m05 vdd b z   vdd p w=1.43u l=0.13u ad=0.360926p pd=2.36167u as=0.3003p   ps=1.885u  
m06 z   b vdd vdd p w=0.99u l=0.13u ad=0.2079p   pd=1.305u   as=0.249872p ps=1.635u  
m07 vdd a z   vdd p w=0.99u l=0.13u ad=0.249872p pd=1.635u   as=0.2079p   ps=1.305u  
m08 w1  a vss vss n w=1.1u  l=0.13u ad=0.14025p  pd=1.355u   as=0.457875p ps=2.4825u 
m09 z   b w1  vss n w=1.1u  l=0.13u ad=0.231p    pd=1.52u    as=0.14025p  ps=1.355u  
m10 w2  b z   vss n w=1.1u  l=0.13u ad=0.14025p  pd=1.355u   as=0.231p    ps=1.52u   
m11 vss a w2  vss n w=1.1u  l=0.13u ad=0.457875p pd=2.4825u  as=0.14025p  ps=1.355u  
m12 w3  a vss vss n w=1.1u  l=0.13u ad=0.14025p  pd=1.355u   as=0.457875p ps=2.4825u 
m13 z   b w3  vss n w=1.1u  l=0.13u ad=0.231p    pd=1.52u    as=0.14025p  ps=1.355u  
m14 w4  b z   vss n w=1.1u  l=0.13u ad=0.14025p  pd=1.355u   as=0.231p    ps=1.52u   
m15 vss a w4  vss n w=1.1u  l=0.13u ad=0.457875p pd=2.4825u  as=0.14025p  ps=1.355u  
C0  a   z   0.378f
C1  b   z   0.221f
C2  a   w1  0.006f
C3  a   w2  0.006f
C4  z   w1  0.009f
C5  a   w3  0.006f
C6  z   w2  0.009f
C7  a   w4  0.006f
C8  z   w3  0.009f
C9  vdd a   0.019f
C10 vdd b   0.037f
C11 vdd z   0.132f
C12 a   b   0.663f
C13 w4  vss 0.010f
C14 w3  vss 0.008f
C15 w2  vss 0.009f
C16 w1  vss 0.009f
C17 z   vss 0.606f
C18 b   vss 0.300f
C19 a   vss 0.391f
.ends
