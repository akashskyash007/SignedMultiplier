.subckt iv1v7x1 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v7x1.ext -        technology: scmos
m00 z   a vdd vdd p w=0.99u  l=0.13u ad=0.29865p pd=2.73u as=0.5709p   ps=4.16u
m01 vss a z   vss n w=0.495u l=0.13u ad=0.41855p pd=3.39u as=0.167475p ps=1.74u
C0 vdd a   0.063f
C1 a   z   0.083f
C2 z   vss 0.114f
C3 a   vss 0.154f
.ends
