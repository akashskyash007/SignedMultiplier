.subckt nr2_x2 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2_x2.ext -        technology: scmos
m00 w1  a vdd vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=1.04033p  ps=5.26u 
m01 z   b w1  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.675u as=0.332475p ps=2.455u
m02 w2  b z   vdd p w=2.145u l=0.13u ad=0.332475p pd=2.455u as=0.568425p ps=2.675u
m03 vdd a w2  vdd p w=2.145u l=0.13u ad=1.04033p  pd=5.26u  as=0.332475p ps=2.455u
m04 z   a vss vss n w=1.155u l=0.13u ad=0.306075p pd=1.685u as=0.560175p ps=3.28u 
m05 vss b z   vss n w=1.155u l=0.13u ad=0.560175p pd=3.28u  as=0.306075p ps=1.685u
C0  z   w3  0.044f
C1  w2  w4  0.005f
C2  a   vdd 0.020f
C3  w1  w5  0.006f
C4  z   w6  0.009f
C5  w2  w3  0.001f
C6  b   vdd 0.020f
C7  z   w5  0.053f
C8  a   z   0.099f
C9  w2  w5  0.006f
C10 vdd w1  0.010f
C11 b   z   0.042f
C12 w4  w5  0.166f
C13 a   w4  0.005f
C14 b   w2  0.017f
C15 vdd z   0.053f
C16 w3  w5  0.166f
C17 a   w3  0.003f
C18 b   w4  0.005f
C19 w1  z   0.012f
C20 vdd w2  0.010f
C21 w6  w5  0.166f
C22 a   w6  0.036f
C23 b   w3  0.012f
C24 vdd w4  0.025f
C25 b   w6  0.001f
C26 vdd w3  0.010f
C27 w1  w4  0.005f
C28 a   w5  0.010f
C29 w1  w3  0.001f
C30 b   w5  0.022f
C31 z   w4  0.008f
C32 a   b   0.303f
C33 vdd w5  0.059f
C34 w5  vss 1.027f
C35 w6  vss 0.179f
C36 w3  vss 0.167f
C37 w4  vss 0.167f
C38 z   vss 0.121f
C40 b   vss 0.096f
C41 a   vss 0.145f
.ends
