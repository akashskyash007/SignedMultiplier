.subckt nd2ab_x1 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nd2ab_x1.ext -        technology: scmos
m00 vdd b  bn  vdd p w=0.99u  l=0.13u ad=0.339726p pd=1.96105u as=0.3168p   ps=2.84u   
m01 z   bn vdd vdd p w=1.1u   l=0.13u ad=0.2915p   pd=1.63u    as=0.377474p ps=2.17895u
m02 vdd an z   vdd p w=1.1u   l=0.13u ad=0.377474p pd=2.17895u as=0.2915p   ps=1.63u   
m03 an  a  vdd vdd p w=0.99u  l=0.13u ad=0.3168p   pd=2.84u    as=0.339726p ps=1.96105u
m04 bn  b  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.21285p  ps=1.48371u
m05 an  a  vss vss n w=0.495u l=0.13u ad=0.185625p pd=1.85u    as=0.21285p  ps=1.48371u
m06 w1  bn z   vss n w=0.935u l=0.13u ad=0.144925p pd=1.245u   as=0.302225p ps=2.73u   
m07 vss an w1  vss n w=0.935u l=0.13u ad=0.40205p  pd=2.80257u as=0.144925p ps=1.245u  
C0  z   w2  0.052f
C1  vdd a   0.057f
C2  a   w2  0.025f
C3  b   z   0.041f
C4  bn  an  0.111f
C5  w1  w2  0.004f
C6  vdd w3  0.021f
C7  bn  z   0.081f
C8  w3  w2  0.166f
C9  vdd w4  0.009f
C10 an  z   0.012f
C11 w4  w2  0.166f
C12 b   w3  0.011f
C13 an  a   0.139f
C14 w5  w2  0.166f
C15 vdd w2  0.038f
C16 b   w4  0.011f
C17 bn  w3  0.001f
C18 z   a   0.067f
C19 b   w5  0.002f
C20 bn  w4  0.011f
C21 an  w3  0.001f
C22 z   w1  0.009f
C23 vdd b   0.092f
C24 b   w2  0.019f
C25 bn  w5  0.011f
C26 an  w4  0.011f
C27 bn  w2  0.022f
C28 an  w5  0.033f
C29 z   w4  0.013f
C30 an  w2  0.020f
C31 z   w5  0.009f
C32 a   w4  0.011f
C33 b   bn  0.075f
C34 w2  vss 1.022f
C35 w5  vss 0.178f
C36 w4  vss 0.165f
C37 w3  vss 0.183f
C38 w1  vss 0.009f
C39 a   vss 0.069f
C40 z   vss 0.117f
C41 an  vss 0.140f
C42 bn  vss 0.124f
C43 b   vss 0.059f
.ends
