.subckt nr2v1x2 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2v1x2.ext -        technology: scmos
m00 w1  a vdd vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u   as=0.611325p ps=3.83u  
m01 z   b w1  vdd p w=1.485u l=0.13u ad=0.31185p  pd=1.905u  as=0.189338p ps=1.74u  
m02 w2  b z   vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u   as=0.31185p  ps=1.905u 
m03 vdd a w2  vdd p w=1.485u l=0.13u ad=0.611325p pd=3.83u   as=0.189338p ps=1.74u  
m04 z   a vss vss n w=0.715u l=0.13u ad=0.160738p pd=1.3275u as=0.218969p ps=1.685u 
m05 vss b z   vss n w=0.715u l=0.13u ad=0.218969p pd=1.685u  as=0.160738p ps=1.3275u
m06 z   b vss vss n w=0.715u l=0.13u ad=0.160738p pd=1.3275u as=0.218969p ps=1.685u 
m07 vss a z   vss n w=0.715u l=0.13u ad=0.218969p pd=1.685u  as=0.160738p ps=1.3275u
C0  vdd a   0.014f
C1  vdd b   0.037f
C2  vdd w1  0.003f
C3  a   b   0.373f
C4  vdd z   0.033f
C5  vdd w2  0.003f
C6  a   z   0.198f
C7  b   z   0.044f
C8  b   w2  0.006f
C9  w1  z   0.009f
C10 w2  vss 0.010f
C11 z   vss 0.349f
C12 w1  vss 0.010f
C13 b   vss 0.175f
C14 a   vss 0.262f
.ends
