.subckt no4_x4 i0 i1 i2 i3 nq vdd vss
*05-JAN-08 SPICE3       file   created      from no4_x4.ext -        technology: scmos
m00 w1  i1 w2  vdd p w=2.19u l=0.13u ad=0.33945p  pd=2.5u     as=1.17055p  ps=5.67u   
m01 w3  i0 w1  vdd p w=2.19u l=0.13u ad=0.33945p  pd=2.5u     as=0.33945p  ps=2.5u    
m02 w4  i2 w3  vdd p w=2.19u l=0.13u ad=0.33945p  pd=2.5u     as=0.33945p  ps=2.5u    
m03 vdd i3 w4  vdd p w=2.19u l=0.13u ad=0.906163p pd=3.36219u as=0.33945p  ps=2.5u    
m04 nq  w5 vdd vdd p w=2.19u l=0.13u ad=0.58035p  pd=2.72u    as=0.906163p ps=3.36219u
m05 vdd w5 nq  vdd p w=2.19u l=0.13u ad=0.906163p pd=3.36219u as=0.58035p  ps=2.72u   
m06 w5  w2 vdd vdd p w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.451012p ps=1.67342u
m07 w2  i1 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.229832p ps=1.41086u
m08 vss i0 w2  vss n w=0.54u l=0.13u ad=0.229832p pd=1.41086u as=0.1431p   ps=1.07u   
m09 w2  i2 vss vss n w=0.54u l=0.13u ad=0.1431p   pd=1.07u    as=0.229832p ps=1.41086u
m10 vss i3 w2  vss n w=0.54u l=0.13u ad=0.229832p pd=1.41086u as=0.1431p   ps=1.07u   
m11 nq  w5 vss vss n w=1.09u l=0.13u ad=0.35925p  pd=2.06u    as=0.46392p  ps=2.84785u
m12 vss w5 nq  vss n w=1.09u l=0.13u ad=0.46392p  pd=2.84785u as=0.35925p  ps=2.06u   
m13 w5  w2 vss vss n w=0.54u l=0.13u ad=0.2295p   pd=1.93u    as=0.229832p ps=1.41086u
C0  i3  w2  0.014f
C1  i0  w3  0.031f
C2  vdd i1  0.021f
C3  w5  w2  0.164f
C4  vdd i0  0.021f
C5  i2  w4  0.052f
C6  vdd i2  0.021f
C7  vdd i3  0.072f
C8  i1  i0  0.261f
C9  vdd w5  0.046f
C10 i1  i2  0.002f
C11 w5  nq  0.020f
C12 vdd w2  0.028f
C13 i0  i2  0.271f
C14 w2  nq  0.076f
C15 vdd w1  0.011f
C16 i1  w2  0.182f
C17 vdd w3  0.011f
C18 i2  i3  0.277f
C19 i0  w2  0.014f
C20 i1  w1  0.019f
C21 vdd w4  0.011f
C22 i2  w2  0.015f
C23 vdd nq  0.076f
C24 i3  w5  0.006f
C25 nq  vss 0.105f
C26 w4  vss 0.007f
C27 w3  vss 0.010f
C28 w1  vss 0.011f
C29 w2  vss 0.444f
C30 w5  vss 0.302f
C31 i3  vss 0.139f
C32 i2  vss 0.129f
C33 i0  vss 0.141f
C34 i1  vss 0.140f
.ends
