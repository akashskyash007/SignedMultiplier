* Spice description of o4_x2
* Spice driver version 134999461
* Date  5/01/2008 at 15:28:54
* sxlib 0.13um values
.subckt o4_x2 i0 i1 i2 i3 q vdd vss
Mtr_00001 sig3  i2    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00002 vss   i3    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00003 vss   i0    sig3  vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00004 sig3  i1    vss   vss n  L=0.12U  W=0.54U  AS=0.1431P   AD=0.1431P   PS=1.61U   PD=1.61U
Mtr_00005 q     sig3  vss   vss n  L=0.12U  W=1.09U  AS=0.28885P  AD=0.28885P  PS=2.71U   PD=2.71U
Mtr_00006 sig6  i3    sig3  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00007 sig7  i1    sig6  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00008 sig5  i0    sig7  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00009 vdd   i2    sig5  vdd p  L=0.12U  W=1.64U  AS=0.4346P   AD=0.4346P   PS=3.81U   PD=3.81U
Mtr_00010 vdd   sig3  q     vdd p  L=0.12U  W=2.19U  AS=0.58035P  AD=0.58035P  PS=4.91U   PD=4.91U
C8  i0    vss   0.882f
C10 i1    vss   0.797f
C9  i2    vss   0.880f
C11 i3    vss   0.746f
C2  q     vss   0.933f
C3  sig3  vss   1.187f
.ends
