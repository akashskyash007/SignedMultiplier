.subckt nmx2_x1 cmd i0 i1 nq vdd vss
*05-JAN-08 SPICE3       file   created      from nmx2_x1.ext -        technology: scmos
m00 vdd cmd w1  vdd p w=1.1u   l=0.13u ad=0.397375p pd=2.14167u as=0.473p    ps=3.06u   
m01 w2  i0  vdd vdd p w=2.09u  l=0.13u ad=0.440393p pd=2.53169u as=0.755013p ps=4.06917u
m02 nq  cmd w2  vdd p w=2.145u l=0.13u ad=0.568425p pd=2.70974u as=0.451982p ps=2.59831u
m03 w3  w1  nq  vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u    as=0.55385p  ps=2.64026u
m04 vdd i1  w3  vdd p w=2.09u  l=0.13u ad=0.755013p pd=4.06917u as=0.55385p  ps=2.62u   
m05 vss cmd w1  vss n w=0.55u  l=0.13u ad=0.199016p pd=1.30217u as=0.2365p   ps=1.96u   
m06 w4  i0  vss vss n w=0.99u  l=0.13u ad=0.2079p   pd=1.41u    as=0.358229p ps=2.34391u
m07 nq  w1  w4  vss n w=0.99u  l=0.13u ad=0.26235p  pd=1.53243u as=0.2079p   ps=1.41u   
m08 w5  cmd nq  vss n w=1.045u l=0.13u ad=0.276925p pd=1.61757u as=0.276925p ps=1.61757u
m09 vss i1  w5  vss n w=0.99u  l=0.13u ad=0.358229p pd=2.34391u as=0.26235p  ps=1.53243u
C0  vdd nq  0.017f
C1  w1  w4  0.015f
C2  vdd w3  0.017f
C3  i0  cmd 0.256f
C4  i0  w1  0.165f
C5  cmd w1  0.139f
C6  i0  vdd 0.044f
C7  cmd i1  0.030f
C8  cmd vdd 0.013f
C9  w1  i1  0.152f
C10 cmd w2  0.035f
C11 w1  vdd 0.154f
C12 cmd nq  0.110f
C13 w1  w2  0.014f
C14 i1  vdd 0.054f
C15 w1  nq  0.139f
C16 i1  nq  0.012f
C17 w1  w3  0.050f
C18 vdd w2  0.014f
C19 w5  vss 0.029f
C20 w4  vss 0.020f
C21 w3  vss 0.019f
C22 nq  vss 0.137f
C23 w2  vss 0.016f
C25 i1  vss 0.163f
C26 w1  vss 0.476f
C27 cmd vss 0.263f
C28 i0  vss 0.126f
.ends
