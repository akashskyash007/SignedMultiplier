.subckt aon21bv0x4 a1 a2 b vdd vss z
*01-JAN-08 SPICE3       file   created      from aon21bv0x4.ext -        technology: scmos
m00 z   an vdd vdd p w=1.43u  l=0.13u ad=0.3003p    pd=1.885u   as=0.405494p  ps=2.691u  
m01 vdd b  z   vdd p w=1.43u  l=0.13u ad=0.405494p  pd=2.691u   as=0.3003p    ps=1.885u  
m02 z   b  vdd vdd p w=1.21u  l=0.13u ad=0.2541p    pd=1.595u   as=0.343111p  ps=2.277u  
m03 vdd an z   vdd p w=1.21u  l=0.13u ad=0.343111p  pd=2.277u   as=0.2541p    ps=1.595u  
m04 an  a1 vdd vdd p w=0.935u l=0.13u ad=0.19635p   pd=1.38125u as=0.265131p  ps=1.7595u 
m05 vdd a2 an  vdd p w=0.935u l=0.13u ad=0.265131p  pd=1.7595u  as=0.19635p   ps=1.38125u
m06 an  a2 vdd vdd p w=0.825u l=0.13u ad=0.17325p   pd=1.21875u as=0.233939p  ps=1.5525u 
m07 vdd a1 an  vdd p w=0.825u l=0.13u ad=0.233939p  pd=1.5525u  as=0.17325p   ps=1.21875u
m08 w1  an vss vss n w=1.1u   l=0.13u ad=0.14025p   pd=1.355u   as=0.513333p  ps=2.87576u
m09 z   b  w1  vss n w=1.1u   l=0.13u ad=0.231p     pd=1.52u    as=0.14025p   ps=1.355u  
m10 w2  b  z   vss n w=1.1u   l=0.13u ad=0.14025p   pd=1.355u   as=0.231p     ps=1.52u   
m11 vss an w2  vss n w=1.1u   l=0.13u ad=0.513333p  pd=2.87576u as=0.14025p   ps=1.355u  
m12 w3  a1 vss vss n w=0.825u l=0.13u ad=0.105188p  pd=1.08u    as=0.385p     ps=2.15682u
m13 an  a2 w3  vss n w=0.825u l=0.13u ad=0.180231p  pd=1.43654u as=0.105188p  ps=1.08u   
m14 w4  a2 an  vss n w=0.605u l=0.13u ad=0.0771375p pd=0.86u    as=0.132169p  ps=1.05346u
m15 vss a1 w4  vss n w=0.605u l=0.13u ad=0.282333p  pd=1.58167u as=0.0771375p ps=0.86u   
C0  vdd z   0.200f
C1  an  a1  0.228f
C2  an  a2  0.057f
C3  an  z   0.164f
C4  an  w1  0.008f
C5  b   z   0.083f
C6  a1  a2  0.283f
C7  an  w2  0.008f
C8  an  w3  0.017f
C9  vdd an  0.150f
C10 z   w1  0.009f
C11 vdd b   0.028f
C12 vdd a1  0.033f
C13 a2  w4  0.010f
C14 vdd a2  0.007f
C15 an  b   0.288f
C16 w4  vss 0.003f
C17 w3  vss 0.004f
C18 w2  vss 0.011f
C19 w1  vss 0.009f
C20 z   vss 0.311f
C21 a2  vss 0.260f
C22 a1  vss 0.200f
C23 b   vss 0.150f
C24 an  vss 0.369f
.ends
