.subckt nr2v0x1 a b vdd vss z
*10-JAN-08 SPICE3       file   created      from nr2v0x1.ext -        technology: scmos
m00 w1  a vdd vdd p w=1.54u l=0.13u ad=0.517p  pd=2.73u as=0.5775p ps=3.83u
m01 z   b w1  vdd p w=1.54u l=0.13u ad=0.5775p pd=3.83u as=0.517p  ps=2.73u
m02 z   a vss vss n w=1.1u  l=0.13u ad=0.4004p pd=2.29u as=0.4125p ps=2.95u
m03 vss b z   vss n w=1.1u  l=0.13u ad=0.4125p pd=2.95u as=0.4004p ps=2.29u
C0  a   b   0.089f
C1  a   z   0.091f
C2  w1  z   0.022f
C3  b   z   0.126f
C4  vdd a   0.038f
C5  vdd w1  0.010f
C6  vdd b   0.007f
C7  z   vss 0.123f
C8  b   vss 0.178f
C9  w1  vss 0.018f
C10 a   vss 0.178f
.ends
