.subckt vfeed2 vdd vss
*10-JAN-08 SPICE3       file   created      from vfeed2.ext -        technology: scmos
m00 w1  vdd w2  vdd p w=1.43u l=0.13u ad=0.37895p pd=1.96u as=0.53625p ps=3.61u
m01 w3  vdd w1  vdd p w=1.43u l=0.13u ad=0.53625p pd=3.61u as=0.37895p ps=1.96u
m02 w4  vdd w5  vdd p w=1.43u l=0.13u ad=0.37895p pd=1.96u as=0.53625p ps=3.61u
m03 w6  vdd w4  vdd p w=1.43u l=0.13u ad=0.53625p pd=3.61u as=0.37895p ps=1.96u
m04 w7  vss w8  vss n w=0.99u l=0.13u ad=0.26235p pd=1.52u as=0.37125p ps=2.73u
m05 w9  vss w7  vss n w=0.99u l=0.13u ad=0.37125p pd=2.73u as=0.26235p ps=1.52u
m06 w10 vss w11 vss n w=0.99u l=0.13u ad=0.26235p pd=1.52u as=0.37125p ps=2.73u
m07 w12 vss w10 vss n w=0.99u l=0.13u ad=0.37125p pd=2.73u as=0.26235p ps=1.52u
C0  w12 vss 0.011f
C1  w10 vss 0.013f
C2  w11 vss 0.011f
C3  w9  vss 0.011f
C4  w7  vss 0.013f
C5  w8  vss 0.011f
C6  w6  vss 0.014f
C7  w4  vss 0.017f
C8  w5  vss 0.014f
C9  w3  vss 0.014f
C10 w1  vss 0.017f
C11 w2  vss 0.014f
.ends
