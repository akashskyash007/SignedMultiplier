.subckt nr3v0x2 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from nr3v0x2.ext -        technology: scmos
m00 w1  c z   vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.365292p ps=2.51u   
m01 w2  b w1  vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.189338p ps=1.74u   
m02 vdd a w2  vdd p w=1.485u l=0.13u ad=0.393525p pd=2.51u    as=0.189338p ps=1.74u   
m03 w3  a vdd vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.393525p ps=2.51u   
m04 w4  b w3  vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.189338p ps=1.74u   
m05 z   c w4  vdd p w=1.485u l=0.13u ad=0.365292p pd=2.51u    as=0.189338p ps=1.74u   
m06 w5  c z   vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.365292p ps=2.51u   
m07 w6  b w5  vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u    as=0.189338p ps=1.74u   
m08 vdd a w6  vdd p w=1.485u l=0.13u ad=0.393525p pd=2.51u    as=0.189338p ps=1.74u   
m09 vss c z   vss n w=0.825u l=0.13u ad=0.23375p  pd=1.66667u as=0.200475p ps=1.63u   
m10 z   b vss vss n w=0.825u l=0.13u ad=0.200475p pd=1.63u    as=0.23375p  ps=1.66667u
m11 vss a z   vss n w=0.825u l=0.13u ad=0.23375p  pd=1.66667u as=0.200475p ps=1.63u   
C0  vdd w4  0.004f
C1  c   w1  0.005f
C2  b   z   0.051f
C3  c   w2  0.005f
C4  a   z   0.013f
C5  c   vdd 0.030f
C6  w5  vdd 0.004f
C7  c   w3  0.005f
C8  z   w1  0.009f
C9  b   vdd 0.021f
C10 c   w4  0.005f
C11 z   w2  0.009f
C12 a   vdd 0.021f
C13 z   vdd 0.064f
C14 z   w3  0.009f
C15 w1  vdd 0.004f
C16 w5  c   0.004f
C17 z   w4  0.009f
C18 w2  vdd 0.004f
C19 c   b   0.355f
C20 c   a   0.243f
C21 vdd w3  0.004f
C22 w6  vdd 0.004f
C23 c   z   0.324f
C24 b   a   0.459f
C25 w5  z   0.005f
C26 w6  vss 0.011f
C27 w5  vss 0.008f
C28 w4  vss 0.007f
C29 w3  vss 0.008f
C31 w2  vss 0.009f
C32 w1  vss 0.007f
C33 z   vss 0.370f
C34 a   vss 0.219f
C35 b   vss 0.339f
C36 c   vss 0.196f
.ends
