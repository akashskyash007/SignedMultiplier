* Spice description of rowend_x0
* Spice driver version 134999461
* Date  5/01/2008 at 15:37:00
* ssxlib 0.13um values
.subckt rowend_x0 vdd vss
.ends
