.subckt aon22_x1 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from aon22_x1.ext -        technology: scmos
m00 z   zn vdd vdd p w=1.1u  l=0.13u ad=0.41855p  pd=3.06u    as=0.435188p ps=2.64167u
m01 zn  b1 n3  vdd p w=1.43u l=0.13u ad=0.37895p  pd=1.96u    as=0.426594p ps=2.84u   
m02 n3  b2 zn  vdd p w=1.43u l=0.13u ad=0.426594p pd=2.84u    as=0.37895p  ps=1.96u   
m03 vdd a2 n3  vdd p w=1.43u l=0.13u ad=0.565744p pd=3.43417u as=0.426594p ps=2.84u   
m04 n3  a1 vdd vdd p w=1.43u l=0.13u ad=0.426594p pd=2.84u    as=0.565744p ps=3.43417u
m05 vss zn z   vss n w=0.55u l=0.13u ad=0.407324p pd=2.02059u as=0.2002p   ps=1.96u   
m06 w1  b1 vss vss n w=0.66u l=0.13u ad=0.1023p   pd=0.97u    as=0.488788p ps=2.42471u
m07 zn  b2 w1  vss n w=0.66u l=0.13u ad=0.1749p   pd=1.19u    as=0.1023p   ps=0.97u   
m08 w2  a2 zn  vss n w=0.66u l=0.13u ad=0.1023p   pd=0.97u    as=0.1749p   ps=1.19u   
m09 vss a1 w2  vss n w=0.66u l=0.13u ad=0.488788p pd=2.42471u as=0.1023p   ps=0.97u   
C0  w3  w4  0.166f
C1  w4  zn  0.068f
C2  w5  z   0.010f
C3  w2  w4  0.005f
C4  w3  vdd 0.011f
C5  b1  a1  0.019f
C6  b2  a2  0.181f
C7  w1  zn  0.010f
C8  w6  w4  0.166f
C9  w4  z   0.026f
C10 w6  vdd 0.007f
C11 vdd z   0.008f
C12 b1  n3  0.007f
C13 b2  a1  0.003f
C14 w5  w4  0.166f
C15 w3  b1  0.001f
C16 b2  n3  0.054f
C17 b1  zn  0.179f
C18 a2  a1  0.192f
C19 w4  vdd 0.052f
C20 w3  b2  0.001f
C21 w6  b1  0.001f
C22 b2  zn  0.051f
C23 a2  n3  0.038f
C24 w1  w4  0.003f
C25 w3  a2  0.001f
C26 w5  b1  0.014f
C27 w6  b2  0.020f
C28 a1  n3  0.007f
C29 w4  b1  0.021f
C30 w3  a1  0.001f
C31 w5  b2  0.013f
C32 w6  a2  0.021f
C33 w2  a1  0.005f
C34 vdd b1  0.002f
C35 w1  b1  0.005f
C36 w4  b2  0.014f
C37 w6  a1  0.001f
C38 w5  a2  0.010f
C39 w3  n3  0.061f
C40 n3  zn  0.069f
C41 vdd b2  0.002f
C42 w4  a2  0.013f
C43 w5  a1  0.012f
C44 w6  n3  0.008f
C45 w3  zn  0.006f
C46 vdd a2  0.041f
C47 w4  a1  0.023f
C48 w6  zn  0.015f
C49 zn  z   0.078f
C50 vdd a1  0.002f
C51 b1  b2  0.178f
C52 w4  n3  0.018f
C53 w5  zn  0.011f
C54 w6  z   0.030f
C55 vdd n3  0.155f
C56 w4  vss 0.985f
C57 w5  vss 0.173f
C58 w6  vss 0.156f
C59 w3  vss 0.160f
C60 z   vss 0.078f
C61 zn  vss 0.248f
C62 n3  vss 0.002f
C63 a1  vss 0.102f
C64 a2  vss 0.081f
C65 b2  vss 0.089f
C66 b1  vss 0.096f
.ends
