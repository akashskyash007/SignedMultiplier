.subckt on12_x1 i0 i1 q vdd vss
*05-JAN-08 SPICE3       file   created      from on12_x1.ext -        technology: scmos
m00 vdd i1 w1  vdd p w=1.09u l=0.13u ad=0.44085p  pd=2.67667u as=0.46325p  ps=3.03u   
m01 q   w1 vdd vdd p w=1.09u l=0.13u ad=0.28885p  pd=1.62u    as=0.44085p  ps=2.67667u
m02 vdd i0 q   vdd p w=1.09u l=0.13u ad=0.44085p  pd=2.67667u as=0.28885p  ps=1.62u   
m03 vss i1 w1  vss n w=0.54u l=0.13u ad=0.218899p pd=1.36491u as=0.2295p   ps=1.93u   
m04 w2  w1 vss vss n w=1.09u l=0.13u ad=0.16895p  pd=1.4u     as=0.441851p ps=2.75509u
m05 q   i0 w2  vss n w=1.09u l=0.13u ad=0.46325p  pd=3.03u    as=0.16895p  ps=1.4u    
C0  vdd i1  0.046f
C1  vdd w1  0.012f
C2  vdd i0  0.046f
C3  i1  w1  0.191f
C4  i1  i0  0.002f
C5  vdd q   0.010f
C6  i1  q   0.166f
C7  w1  i0  0.096f
C8  i0  q   0.180f
C9  q   w2  0.020f
C10 w2  vss 0.006f
C11 q   vss 0.131f
C12 i0  vss 0.152f
C13 w1  vss 0.235f
C14 i1  vss 0.203f
.ends
