.subckt nr2_x05 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from nr2_x05.ext -        technology: scmos
m00 w1  b z   vdd p w=1.21u l=0.13u ad=0.18755p pd=1.52u as=0.4477p  ps=3.28u
m01 vdd a w1  vdd p w=1.21u l=0.13u ad=0.58685p pd=3.39u as=0.18755p ps=1.52u
m02 z   b vss vss n w=0.33u l=0.13u ad=0.08745p pd=0.86u as=0.1419p  ps=1.52u
m03 vss a z   vss n w=0.33u l=0.13u ad=0.1419p  pd=1.52u as=0.08745p ps=0.86u
C0 vdd a   0.031f
C1 b   a   0.172f
C2 b   z   0.071f
C3 a   z   0.041f
C4 a   w1  0.015f
C5 w1  vss 0.007f
C6 z   vss 0.147f
C7 a   vss 0.115f
C8 b   vss 0.160f
.ends
