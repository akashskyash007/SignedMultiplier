.subckt vfeed4 vdd vss
*04-JAN-08 SPICE3       file   created      from vfeed4.ext -        technology: scmos
.ends
