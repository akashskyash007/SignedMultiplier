.subckt nr2v0x3 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from nr2v0x3.ext -        technology: scmos
m00 w1  b z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.37785p   ps=2.58333u 
m01 vdd a w1  vdd p w=1.54u  l=0.13u ad=0.436333p pd=2.62u    as=0.19635p   ps=1.795u   
m02 w2  a vdd vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.436333p  ps=2.62u    
m03 z   b w2  vdd p w=1.54u  l=0.13u ad=0.37785p  pd=2.58333u as=0.19635p   ps=1.795u   
m04 w3  b z   vdd p w=1.54u  l=0.13u ad=0.19635p  pd=1.795u   as=0.37785p   ps=2.58333u 
m05 vdd a w3  vdd p w=1.54u  l=0.13u ad=0.436333p pd=2.62u    as=0.19635p   ps=1.795u   
m06 z   b vss vss n w=0.715u l=0.13u ad=0.156704p pd=1.28917u as=0.306631p  ps=2.12333u 
m07 vss a z   vss n w=0.935u l=0.13u ad=0.400979p pd=2.77667u as=0.204921p  ps=1.68583u 
m08 z   b vss vss n w=0.605u l=0.13u ad=0.132596p pd=1.09083u as=0.259457p  ps=1.79667u 
m09 vss a z   vss n w=0.385u l=0.13u ad=0.165109p pd=1.14333u as=0.0843792p ps=0.694167u
C0  vdd w2  0.004f
C1  vdd w3  0.004f
C2  b   a   0.401f
C3  b   z   0.173f
C4  a   z   0.104f
C5  b   vdd 0.021f
C6  z   w1  0.009f
C7  a   vdd 0.034f
C8  a   w2  0.006f
C9  z   vdd 0.058f
C10 a   w3  0.006f
C11 z   w2  0.009f
C12 w1  vdd 0.004f
C13 w3  vss 0.008f
C14 w2  vss 0.007f
C16 w1  vss 0.008f
C17 z   vss 0.391f
C18 a   vss 0.215f
C19 b   vss 0.204f
.ends
