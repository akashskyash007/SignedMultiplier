.subckt an2_x1 a b vdd vss z
*04-JAN-08 SPICE3       file   created      from an2_x1.ext -        technology: scmos
m00 vdd zn z   vdd p w=1.1u  l=0.13u ad=0.459039p pd=2.85385u as=0.41855p  ps=3.06u   
m01 zn  a  vdd vdd p w=0.88u l=0.13u ad=0.2332p   pd=1.41u    as=0.367231p ps=2.28308u
m02 vdd b  zn  vdd p w=0.88u l=0.13u ad=0.367231p pd=2.28308u as=0.2332p   ps=1.41u   
m03 vss zn z   vss n w=0.55u l=0.13u ad=0.26675p  pd=1.49583u as=0.2002p   ps=1.96u   
m04 w1  a  vss vss n w=0.77u l=0.13u ad=0.11935p  pd=1.08u    as=0.37345p  ps=2.09417u
m05 zn  b  w1  vss n w=0.77u l=0.13u ad=0.3311p   pd=2.4u     as=0.11935p  ps=1.08u   
C0  vdd w2  0.034f
C1  z   w3  0.001f
C2  zn  w4  0.031f
C3  zn  w5  0.013f
C4  z   w4  0.013f
C5  zn  w2  0.035f
C6  z   w5  0.010f
C7  vdd zn  0.015f
C8  z   w2  0.022f
C9  a   w5  0.025f
C10 b   w4  0.010f
C11 vdd z   0.029f
C12 a   w2  0.013f
C13 b   w2  0.018f
C14 vdd b   0.018f
C15 zn  z   0.109f
C16 w1  w2  0.006f
C17 zn  a   0.150f
C18 w3  w2  0.166f
C19 vdd w3  0.021f
C20 zn  b   0.077f
C21 w4  w2  0.166f
C22 vdd w4  0.005f
C23 z   b   0.016f
C24 zn  w1  0.010f
C25 w5  w2  0.166f
C26 zn  w3  0.002f
C27 a   b   0.146f
C28 w2  vss 1.033f
C29 w5  vss 0.181f
C30 w4  vss 0.175f
C31 w3  vss 0.185f
C32 b   vss 0.069f
C33 a   vss 0.087f
C34 z   vss 0.022f
C35 zn  vss 0.157f
.ends
