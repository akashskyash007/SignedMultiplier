.subckt iv1v1x4 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v1x4.ext -        technology: scmos
m00 z   a vdd vdd p w=1.54u  l=0.13u ad=0.3234p   pd=1.96u  as=0.61985p  ps=3.885u
m01 vdd a z   vdd p w=1.54u  l=0.13u ad=0.61985p  pd=3.885u as=0.3234p   ps=1.96u 
m02 z   a vss vss n w=1.045u l=0.13u ad=0.21945p  pd=1.465u as=0.420613p ps=2.895u
m03 vss a z   vss n w=1.045u l=0.13u ad=0.420613p pd=2.895u as=0.21945p  ps=1.465u
C0 vdd a   0.024f
C1 vdd z   0.089f
C2 a   z   0.058f
C3 z   vss 0.241f
C4 a   vss 0.166f
.ends
