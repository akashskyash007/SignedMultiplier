.subckt nd3v0x1 a b c vdd vss z
*01-JAN-08 SPICE3       file   created      from nd3v0x1.ext -        technology: scmos
m00 vdd c z   vdd p w=1.1u l=0.13u ad=0.2915p   pd=1.99667u as=0.277383p ps=1.99667u
m01 z   b vdd vdd p w=1.1u l=0.13u ad=0.277383p pd=1.99667u as=0.2915p   ps=1.99667u
m02 vdd a z   vdd p w=1.1u l=0.13u ad=0.2915p   pd=1.99667u as=0.277383p ps=1.99667u
m03 w1  c z   vss n w=1.1u l=0.13u ad=0.14025p  pd=1.355u   as=0.3278p   ps=2.95u   
m04 w2  b w1  vss n w=1.1u l=0.13u ad=0.14025p  pd=1.355u   as=0.14025p  ps=1.355u  
m05 vss a w2  vss n w=1.1u l=0.13u ad=0.5093p   pd=3.28u    as=0.14025p  ps=1.355u  
C0  vdd c   0.007f
C1  vdd b   0.034f
C2  vdd a   0.007f
C3  vdd z   0.111f
C4  c   b   0.124f
C5  c   a   0.037f
C6  c   z   0.076f
C7  b   a   0.177f
C8  c   w1  0.007f
C9  b   z   0.049f
C10 c   w2  0.005f
C11 w2  vss 0.011f
C12 w1  vss 0.010f
C13 z   vss 0.249f
C14 a   vss 0.152f
C15 b   vss 0.104f
C16 c   vss 0.091f
.ends
