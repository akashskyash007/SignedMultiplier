* Spice description of oai22v0x05
* Spice driver version 134999461
* Date  1/01/2008 at 16:59:05
* vsclib 0.13um values
.subckt oai22v0x05 a1 a2 b1 b2 vdd vss z
M01 vdd   a1    03    vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M02 sig1  a1    vss   vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M03 03    a2    z     vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M04 vss   a2    sig1  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M05 z     b2    sig8  vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M06 sig1  b2    z     vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
M07 sig8  b1    vdd   vdd p  L=0.12U  W=0.88U  AS=0.2332P   AD=0.2332P   PS=2.29U   PD=2.29U
M08 z     b1    sig1  vss n  L=0.12U  W=0.385U AS=0.102025P AD=0.102025P PS=1.3U    PD=1.3U
C7  a1    vss   0.680f
C6  a2    vss   0.566f
C4  b1    vss   0.605f
C5  b2    vss   0.539f
C1  sig1  vss   0.324f
C2  z     vss   0.797f
.ends
