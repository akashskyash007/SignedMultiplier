* Spice description of an3_x2
* Spice driver version 134999461
* Date  4/01/2008 at 18:48:59
* vsxlib 0.13um values
.subckt an3_x2 a b c vdd vss z
M1a 2z    a     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1b vdd   b     2z    vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1c 2z    c     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M1z vdd   2z    z     vdd p  L=0.12U  W=2.09U  AS=0.55385P  AD=0.55385P  PS=4.71U   PD=4.71U
M2a vss   a     sig4  vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2b sig4  b     n2    vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2c n2    c     2z    vss n  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M2z z     2z    vss   vss n  L=0.12U  W=1.045U AS=0.276925P AD=0.276925P PS=2.62U   PD=2.62U
C3  2z    vss   1.240f
C8  a     vss   0.817f
C7  b     vss   0.783f
C6  c     vss   0.881f
C1  z     vss   0.796f
.ends
