.subckt zero_x0 nq vdd vss
*05-JAN-08 SPICE3       file   created      from zero_x0.ext -        technology: scmos
m00 nq vdd vss vss n w=0.55u l=0.13u ad=0.2365p pd=1.96u as=0.297p ps=2.18u
C0 vdd nq  0.132f
C1 nq  vss 0.150f
.ends
