.subckt iv1v1x05 a vdd vss z
*01-JAN-08 SPICE3       file   created      from iv1v1x05.ext -        technology: scmos
m00 z   a vdd vdd p w=0.66u l=0.13u ad=0.2112p pd=2.07u as=0.559075p ps=4.27u
m01 vss a z   vss n w=0.44u l=0.13u ad=0.165p  pd=1.63u as=0.1529p   ps=1.63u
C0 vdd a   0.060f
C1 a   z   0.031f
C2 z   vss 0.101f
C3 a   vss 0.108f
.ends
