* Spice description of an12_x1
* Spice driver version 134999461
* Date  5/01/2008 at 15:01:20
* ssxlib 0.13um values
.subckt an12_x1 i0 i1 q vdd vss
Mtr_00001 vss   i1    sig4  vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00002 q     sig4  vss   vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00003 vss   i0    q     vss n  L=0.12U  W=0.55U  AS=0.14575P  AD=0.14575P  PS=1.63U   PD=1.63U
Mtr_00004 sig4  i1    vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
Mtr_00005 vdd   sig4  sig7  vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
Mtr_00006 sig7  i0    q     vdd p  L=0.12U  W=2.145U AS=0.568425P AD=0.568425P PS=4.82U   PD=4.82U
C3  i0    vss   0.977f
C5  i1    vss   1.081f
C2  q     vss   0.912f
C4  sig4  vss   0.783f
.ends
