* functionality check of iv1v0x4, 0.13um, Berkeley generic bsim3 params
* iv1v0x4_func.cir 2008-01-11:21h03 graham
*
.include ../../../magic/subckt/vgalib013/spice_model.lib
.include ../../../magic/subckt/vgalib013/iv1v0x4.spi
.include ../../../magic/subckt/vgalib013/params.inc
*
x01 va   vdd vss x01z iv1v0x4
x02 va   vdd vss x02z iv1v0x4
*
.param unitcap=1.5f
cx01z  x01z  0 '4*unitcap'
cx02z  x02z  0 '130*4*unitcap'
* 
vdd vdd 0 'vdd'
vss 0 vss 'vss'
vstrobe strobe 0 dc 0 pulse (0 1 '0.97*tPER' '0.01*tPER' '0.01*tPER' '0.01*tPER' 'tPER')
*           00   10     11     01     00     01     11     10     00
*            0    1      0      1      0      1      0      1      0
*                thh_AZ thl_BZ tlh_AZ tll_BZ thh_BZ thl_AZ tlh_BZ tll_AZ
*                 0      1      2      3      4      5      6      7      8
Va  va 0 pwl(0 'vss' 'tRISE'  'vdd' '1*tPER' 'vdd'  '1*tPER+tFALL' 'vss'
+           '2*tPER' 'vss' '2*tPER+tRISE' 'vdd' '3*tPER' 'vdd' '3*tPER+tFALL' 'vss' )

.control
  set width=120 height=500 numdgt=3 noprintscale nobreak noaskquit=1
  tran $tstep 20000p
  linearize
  let a = va / $vdd
  let pa = va + $vdd + 0.3
  let pz = $vdd * (not a) - $vdd - 0.3
* check output is within 10mV of ideal at strobe point
  let perr =  vecmax ( pos ( abs (( pz - x02z + $vdd + 0.3 ) * strobe ) - 0.01 ))
*  plot v(pa) v(pz) v(x01z) v(x02z)
*  print col v(va) v(x01z) v(x02z) > iv1v0x4_func.spo
  if perr > 0
    echo #Error: Functional simulation iv1v0x4_func.cir failed
    echo #Error: Functional simulation iv1v0x4_func.cir failed >> iv1v0x4_func.error
  else
    echo Functional simulation OK
  end
  destroy all
.endc
.end
