.subckt xaon22_x1 a1 a2 b1 b2 vdd vss z
*04-JAN-08 SPICE3       file   created      from xaon22_x1.ext -        technology: scmos
m00 vdd a1 an  vdd p w=1.925u l=0.13u ad=0.721875p pd=2.675u   as=0.552475p ps=3.20667u
m01 an  a2 vdd vdd p w=1.925u l=0.13u ad=0.552475p pd=3.20667u as=0.721875p ps=2.675u  
m02 z   bn an  vdd p w=1.925u l=0.13u ad=0.510125p pd=2.455u   as=0.552475p ps=3.20667u
m03 bn  an z   vdd p w=1.925u l=0.13u ad=0.693642p pd=3.35333u as=0.510125p ps=2.455u  
m04 vdd b1 bn  vdd p w=1.925u l=0.13u ad=0.721875p pd=2.675u   as=0.693642p ps=3.35333u
m05 bn  b2 vdd vdd p w=1.925u l=0.13u ad=0.693642p pd=3.35333u as=0.721875p ps=2.675u  
m06 w1  a1 vss vss n w=1.815u l=0.13u ad=0.281325p pd=2.125u   as=0.679276p ps=3.6523u 
m07 an  a2 w1  vss n w=1.815u l=0.13u ad=0.480975p pd=2.76375u as=0.281325p ps=2.125u  
m08 w2  b2 an  vss n w=1.265u l=0.13u ad=0.196075p pd=1.575u   as=0.335225p ps=1.92625u
m09 z   b1 w2  vss n w=1.265u l=0.13u ad=0.335225p pd=2.0139u  as=0.196075p ps=1.575u  
m10 w3  bn z   vss n w=0.99u  l=0.13u ad=0.15345p  pd=1.3u     as=0.26235p  ps=1.5761u 
m11 vss an w3  vss n w=0.99u  l=0.13u ad=0.370514p pd=1.99216u as=0.15345p  ps=1.3u    
m12 w4  b1 vss vss n w=1.265u l=0.13u ad=0.196075p pd=1.575u   as=0.473435p ps=2.54554u
m13 bn  b2 w4  vss n w=1.265u l=0.13u ad=0.389675p pd=3.39u    as=0.196075p ps=1.575u  
C0  a2  vdd 0.024f
C1  bn  b2  0.048f
C2  an  b1  0.046f
C3  a2  z   0.067f
C4  bn  vdd 0.169f
C5  an  b2  0.016f
C6  bn  z   0.029f
C7  an  vdd 0.180f
C8  b1  b2  0.278f
C9  w2  z   0.015f
C10 w3  an  0.020f
C11 an  z   0.294f
C12 b1  vdd 0.060f
C13 b1  z   0.008f
C14 b2  vdd 0.010f
C15 a1  a2  0.161f
C16 b2  z   0.016f
C17 w4  b2  0.026f
C18 vdd z   0.017f
C19 a2  bn  0.057f
C20 a1  an  0.007f
C21 a2  an  0.092f
C22 bn  an  0.349f
C23 w2  an  0.010f
C24 a2  b2  0.028f
C25 bn  b1  0.168f
C26 a1  vdd 0.010f
C27 w1  vss 0.010f
C28 z   vss 0.017f
C30 b2  vss 0.323f
C31 b1  vss 0.169f
C32 an  vss 0.205f
C33 bn  vss 0.133f
C34 a2  vss 0.082f
C35 a1  vss 0.111f
.ends
