* Spice description of iv1v4x1
* Spice driver version 134999461
* Date  1/01/2008 at 16:45:34
* wsclib 0.13um values
.subckt iv1v4x1 a vdd vss z
M01 z     a     vdd   vdd p  L=0.12U  W=1.32U  AS=0.3498P   AD=0.3498P   PS=3.17U   PD=3.17U
M02 vss   a     z     vss n  L=0.12U  W=0.33U  AS=0.08745P  AD=0.08745P  PS=1.19U   PD=1.19U
C3  a     vss   0.475f
C2  z     vss   0.600f
.ends
