.subckt bf1v0x2 a vdd vss z
*01-JAN-08 SPICE3       file   created      from bf1v0x2.ext -        technology: scmos
m00 vdd an z   vdd p w=1.54u  l=0.13u ad=0.504093p pd=2.78133u as=0.48675p  ps=3.83u   
m01 an  a  vdd vdd p w=0.935u l=0.13u ad=0.284075p pd=2.62u    as=0.306057p ps=1.68867u
m02 vss an z   vss n w=0.77u  l=0.13u ad=0.225225p pd=1.51667u as=0.28875p  ps=2.29u   
m03 an  a  vss vss n w=0.55u  l=0.13u ad=0.18205p  pd=1.85u    as=0.160875p ps=1.08333u
C0 vdd an  0.031f
C1 vdd z   0.055f
C2 an  z   0.136f
C3 an  a   0.156f
C4 a   vss 0.101f
C5 z   vss 0.195f
C6 an  vss 0.140f
.ends
