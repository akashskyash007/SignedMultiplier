.subckt iv1_x4 a vdd vss z
*04-JAN-08 SPICE3       file   created      from iv1_x4.ext -        technology: scmos
m00 z   a vdd vdd p w=2.09u  l=0.13u ad=0.55385p  pd=2.62u  as=1.01365p  ps=5.15u 
m01 vdd a z   vdd p w=2.09u  l=0.13u ad=1.01365p  pd=5.15u  as=0.55385p  ps=2.62u 
m02 z   a vss vss n w=1.045u l=0.13u ad=0.276925p pd=1.575u as=0.506825p ps=3.06u 
m03 vss a z   vss n w=1.045u l=0.13u ad=0.506825p pd=3.06u  as=0.276925p ps=1.575u
C0  z   w1  0.035f
C1  w2  w1  0.166f
C2  w3  w1  0.166f
C3  w4  w1  0.166f
C4  a   vdd 0.043f
C5  a   z   0.092f
C6  vdd z   0.062f
C7  a   w2  0.005f
C8  vdd w2  0.025f
C9  a   w3  0.011f
C10 a   w4  0.011f
C11 vdd w3  0.007f
C12 z   w2  0.008f
C13 a   w1  0.021f
C14 z   w3  0.033f
C15 vdd w1  0.050f
C16 z   w4  0.030f
C17 w1  vss 1.059f
C18 w4  vss 0.184f
C19 w3  vss 0.177f
C20 w2  vss 0.177f
C21 z   vss 0.114f
C23 a   vss 0.138f
.ends
