.subckt xor2v5x1 a b vdd vss z
*01-JAN-08 SPICE3       file   created      from xor2v5x1.ext -        technology: scmos
m00 vdd a  an  vdd p w=0.605u l=0.13u ad=0.222935p pd=1.21434u  as=0.196625p ps=1.96u    
m01 w1  a  vdd vdd p w=1.485u l=0.13u ad=0.189338p pd=1.74u     as=0.547203p ps=2.98066u 
m02 z   bn w1  vdd p w=1.485u l=0.13u ad=0.31185p  pd=1.905u    as=0.189338p ps=1.74u    
m03 w2  an z   vdd p w=1.485u l=0.13u ad=0.31185p  pd=1.905u    as=0.31185p  ps=1.905u   
m04 vdd b  w2  vdd p w=1.485u l=0.13u ad=0.547203p pd=2.98066u  as=0.31185p  ps=1.905u   
m05 bn  b  vdd vdd p w=0.605u l=0.13u ad=0.196625p pd=1.96u     as=0.222935p ps=1.21434u 
m06 vss a  an  vss n w=0.33u  l=0.13u ad=0.08745p  pd=0.738333u as=0.12375p  ps=1.41u    
m07 w3  a  vss vss n w=0.66u  l=0.13u ad=0.08415p  pd=0.915u    as=0.1749p   ps=1.47667u 
m08 z   b  w3  vss n w=0.66u  l=0.13u ad=0.1386p   pd=1.08u     as=0.08415p  ps=0.915u   
m09 w4  bn z   vss n w=0.66u  l=0.13u ad=0.08415p  pd=0.915u    as=0.1386p   ps=1.08u    
m10 vss an w4  vss n w=0.66u  l=0.13u ad=0.1749p   pd=1.47667u  as=0.08415p  ps=0.915u   
m11 bn  b  vss vss n w=0.33u  l=0.13u ad=0.12375p  pd=1.41u     as=0.08745p  ps=0.738333u
C0  b   z   0.024f
C1  an  w2  0.024f
C2  vdd a   0.044f
C3  bn  w4  0.005f
C4  w1  z   0.005f
C5  vdd bn  0.012f
C6  vdd an  0.052f
C7  vdd b   0.007f
C8  a   bn  0.080f
C9  a   an  0.070f
C10 vdd w1  0.004f
C11 vdd z   0.007f
C12 a   b   0.048f
C13 bn  an  0.175f
C14 vdd w2  0.007f
C15 bn  b   0.112f
C16 a   z   0.011f
C17 an  b   0.077f
C18 bn  z   0.087f
C19 an  w1  0.008f
C20 an  z   0.096f
C21 w4  vss 0.004f
C22 w3  vss 0.005f
C23 w2  vss 0.013f
C24 z   vss 0.102f
C25 w1  vss 0.007f
C26 b   vss 0.314f
C27 an  vss 0.221f
C28 bn  vss 0.140f
C29 a   vss 0.175f
.ends
