* Spice description of tie_x0
* Spice driver version 134999461
* Date  4/01/2008 at 19:49:44
* vxlib 0.13um values
.subckt tie_x0 vdd vss
.ends
