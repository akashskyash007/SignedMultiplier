* Spice description of nd2_x1
* Spice driver version 134999461
* Date  4/01/2008 at 19:03:20
* vxlib 0.13um values
.subckt nd2_x1 a b vdd vss z
M1  z     b     vdd   vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M2  vdd   a     z     vdd p  L=0.12U  W=1.1U   AS=0.2915P   AD=0.2915P   PS=2.73U   PD=2.73U
M3  z     b     n1    vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
M4  n1    a     vss   vss n  L=0.12U  W=0.935U AS=0.247775P AD=0.247775P PS=2.4U    PD=2.4U
C5  a     vss   0.740f
C6  b     vss   0.733f
C2  z     vss   0.725f
.ends
